// streaming permutation network
// for degree: 2^16-1
// data parallelism: 256
// data width: 54                                                                                     
 
module switch_2_2(
inData_0,
inData_1,
outData_0,
outData_1,
ctrl,                            
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input ctrl, clk, rst;                   
  input [DATA_WIDTH-1:0] inData_0,
      inData_1;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1;
  
  wire [DATA_WIDTH-1:0] wireIn [1:0];              
  wire [DATA_WIDTH-1:0] wireOut [1:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  
  assign wireOut[0] = (!ctrl) ? wireIn[0] : wireIn[1];    
  assign wireOut[1] = (!ctrl) ? wireIn[1] : wireIn[0];    
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  
endmodule                        


module  counter_512(
in_start,                         
counter_out,                         
clk,                             
rst                              
);                               
  input in_start, clk, rst;                   
  output [8:0] counter_out;            
  
  reg [8:0] counter_r;        
  reg status_couting;        

  assign counter_out = counter_r;        
  
  always@(posedge clk)             
  begin                            
    if(rst) begin                    
      counter_r <= 9'b0;    
      status_couting <= 1'b0;            
    end
    else begin                        
      if (status_couting == 1'b1)                
        counter_r <= counter_r + 1'b1;                   
      if (counter_r[8:0] == 511) begin  
        status_couting <= 1'b0;                 
        counter_r <= 9'b0;         
      end                                    
      if (in_start) begin                     
        status_couting <= 1'b1;                 
      counter_r <= 9'b0;                
      end                                    
    end
  end                              

endmodule                        


module  block_ram_sp(
wen,                              
en,                              
clk,                             
addr,                            
din,                            
dout                             
);                               
  parameter DATA_WIDTH = 54;                                
  parameter ADDR_WIDTH = 8;                                
  parameter RAM_SIZE = 1 << ADDR_WIDTH;                                
  input wen, clk;                   
  input en;                              
  input [ADDR_WIDTH-1:0] addr;                        
  input [DATA_WIDTH-1:0] din;                        
  output reg [DATA_WIDTH-1:0] dout;        
  
  reg [DATA_WIDTH-1:0] ram[RAM_SIZE-1:0];        
  
  always@(posedge clk)             
  begin                            
    // synthesis attribute ram_style of ram is "block" 
  if(en) begin                    
      if(wen)                         
        ram[addr] <= din ;              
      dout <= ram[addr];              
  end
  end                             
  
endmodule                        


module  dist_ram_sp(
wen,                              
clk,                             
addr,                            
din,                            
dout                             
);                               
  parameter DATA_WIDTH = 54;                                
  parameter ADDR_WIDTH = 8;                                
  parameter RAM_SIZE = 1 << ADDR_WIDTH;                                
  input wen, clk;                   
  input [ADDR_WIDTH-1:0] addr;                        
  input [DATA_WIDTH-1:0] din;                        
  output [DATA_WIDTH-1:0] dout;        
  
  reg [DATA_WIDTH-1:0] ram[RAM_SIZE-1:0];        
  
  always@(posedge clk)             
  begin                            
    // synthesis attribute ram_style of ram is "distributed" 
  if(wen)                         
      ram[addr] <= din ;              
  end                             
 
  assign dout = ram[addr];         
  
endmodule                        


module  block_ram_dp(
wen,                              
en,                              
clk,                             
addr_r,                            
addr_w,                            
din,                            
dout                             
);                               
  parameter DATA_WIDTH = 54;                                
  parameter ADDR_WIDTH = 8;                                
  parameter RAM_SIZE = 1 << ADDR_WIDTH;                                
  input wen, clk;                   
  input en;                              
  input [ADDR_WIDTH-1:0] addr_r;                        
  input [ADDR_WIDTH-1:0] addr_w;                        
  input [DATA_WIDTH-1:0] din;                        
  output reg [DATA_WIDTH-1:0] dout;        
  
  reg [DATA_WIDTH-1:0] ram[RAM_SIZE-1:0];        
  
  always@(posedge clk)             
  begin                            
    // synthesis attribute ram_style of ram is "block" 
  if(en) begin                    
      if(wen)                         
        ram[addr_w] <= din ;              
      dout <= ram[addr_r];              
  end
  end                             
  
endmodule                        


module  dist_ram_dp(
wen,                              
clk,                             
addr_r,                            
addr_w,                            
din,                            
dout                             
);                               
  parameter DATA_WIDTH = 54;                                
  parameter ADDR_WIDTH = 8;                                
  parameter RAM_SIZE = 1 << ADDR_WIDTH;                                
  input wen, clk;                   
  input [ADDR_WIDTH-1:0] addr_r;                        
  input [ADDR_WIDTH-1:0] addr_w;                        
  input [DATA_WIDTH-1:0] din;                        
  output [DATA_WIDTH-1:0] dout;        
  
  reg [DATA_WIDTH-1:0] ram[RAM_SIZE-1:0];        
  
  always@(posedge clk)             
  begin                            
    // synthesis attribute ram_style of ram is "distributed" 
  if(wen)                         
      ram[addr_w] <= din ;              
  end                             
 
  assign dout = ram[addr_r];         
  
endmodule                        


module switches_stage_st0_0_L(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
ctrl,                            
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;                   
  input [128-1:0] ctrl;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  switch_2_2 switch_inst_0(.inData_0(wireIn[0]), .inData_1(wireIn[1]), .outData_0(wireOut[0]), .outData_1(wireOut[1]), .ctrl(ctrl[0]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_1(.inData_0(wireIn[2]), .inData_1(wireIn[3]), .outData_0(wireOut[2]), .outData_1(wireOut[3]), .ctrl(ctrl[1]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_2(.inData_0(wireIn[4]), .inData_1(wireIn[5]), .outData_0(wireOut[4]), .outData_1(wireOut[5]), .ctrl(ctrl[2]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_3(.inData_0(wireIn[6]), .inData_1(wireIn[7]), .outData_0(wireOut[6]), .outData_1(wireOut[7]), .ctrl(ctrl[3]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_4(.inData_0(wireIn[8]), .inData_1(wireIn[9]), .outData_0(wireOut[8]), .outData_1(wireOut[9]), .ctrl(ctrl[4]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_5(.inData_0(wireIn[10]), .inData_1(wireIn[11]), .outData_0(wireOut[10]), .outData_1(wireOut[11]), .ctrl(ctrl[5]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_6(.inData_0(wireIn[12]), .inData_1(wireIn[13]), .outData_0(wireOut[12]), .outData_1(wireOut[13]), .ctrl(ctrl[6]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_7(.inData_0(wireIn[14]), .inData_1(wireIn[15]), .outData_0(wireOut[14]), .outData_1(wireOut[15]), .ctrl(ctrl[7]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_8(.inData_0(wireIn[16]), .inData_1(wireIn[17]), .outData_0(wireOut[16]), .outData_1(wireOut[17]), .ctrl(ctrl[8]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_9(.inData_0(wireIn[18]), .inData_1(wireIn[19]), .outData_0(wireOut[18]), .outData_1(wireOut[19]), .ctrl(ctrl[9]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_10(.inData_0(wireIn[20]), .inData_1(wireIn[21]), .outData_0(wireOut[20]), .outData_1(wireOut[21]), .ctrl(ctrl[10]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_11(.inData_0(wireIn[22]), .inData_1(wireIn[23]), .outData_0(wireOut[22]), .outData_1(wireOut[23]), .ctrl(ctrl[11]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_12(.inData_0(wireIn[24]), .inData_1(wireIn[25]), .outData_0(wireOut[24]), .outData_1(wireOut[25]), .ctrl(ctrl[12]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_13(.inData_0(wireIn[26]), .inData_1(wireIn[27]), .outData_0(wireOut[26]), .outData_1(wireOut[27]), .ctrl(ctrl[13]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_14(.inData_0(wireIn[28]), .inData_1(wireIn[29]), .outData_0(wireOut[28]), .outData_1(wireOut[29]), .ctrl(ctrl[14]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_15(.inData_0(wireIn[30]), .inData_1(wireIn[31]), .outData_0(wireOut[30]), .outData_1(wireOut[31]), .ctrl(ctrl[15]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_16(.inData_0(wireIn[32]), .inData_1(wireIn[33]), .outData_0(wireOut[32]), .outData_1(wireOut[33]), .ctrl(ctrl[16]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_17(.inData_0(wireIn[34]), .inData_1(wireIn[35]), .outData_0(wireOut[34]), .outData_1(wireOut[35]), .ctrl(ctrl[17]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_18(.inData_0(wireIn[36]), .inData_1(wireIn[37]), .outData_0(wireOut[36]), .outData_1(wireOut[37]), .ctrl(ctrl[18]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_19(.inData_0(wireIn[38]), .inData_1(wireIn[39]), .outData_0(wireOut[38]), .outData_1(wireOut[39]), .ctrl(ctrl[19]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_20(.inData_0(wireIn[40]), .inData_1(wireIn[41]), .outData_0(wireOut[40]), .outData_1(wireOut[41]), .ctrl(ctrl[20]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_21(.inData_0(wireIn[42]), .inData_1(wireIn[43]), .outData_0(wireOut[42]), .outData_1(wireOut[43]), .ctrl(ctrl[21]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_22(.inData_0(wireIn[44]), .inData_1(wireIn[45]), .outData_0(wireOut[44]), .outData_1(wireOut[45]), .ctrl(ctrl[22]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_23(.inData_0(wireIn[46]), .inData_1(wireIn[47]), .outData_0(wireOut[46]), .outData_1(wireOut[47]), .ctrl(ctrl[23]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_24(.inData_0(wireIn[48]), .inData_1(wireIn[49]), .outData_0(wireOut[48]), .outData_1(wireOut[49]), .ctrl(ctrl[24]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_25(.inData_0(wireIn[50]), .inData_1(wireIn[51]), .outData_0(wireOut[50]), .outData_1(wireOut[51]), .ctrl(ctrl[25]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_26(.inData_0(wireIn[52]), .inData_1(wireIn[53]), .outData_0(wireOut[52]), .outData_1(wireOut[53]), .ctrl(ctrl[26]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_27(.inData_0(wireIn[54]), .inData_1(wireIn[55]), .outData_0(wireOut[54]), .outData_1(wireOut[55]), .ctrl(ctrl[27]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_28(.inData_0(wireIn[56]), .inData_1(wireIn[57]), .outData_0(wireOut[56]), .outData_1(wireOut[57]), .ctrl(ctrl[28]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_29(.inData_0(wireIn[58]), .inData_1(wireIn[59]), .outData_0(wireOut[58]), .outData_1(wireOut[59]), .ctrl(ctrl[29]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_30(.inData_0(wireIn[60]), .inData_1(wireIn[61]), .outData_0(wireOut[60]), .outData_1(wireOut[61]), .ctrl(ctrl[30]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_31(.inData_0(wireIn[62]), .inData_1(wireIn[63]), .outData_0(wireOut[62]), .outData_1(wireOut[63]), .ctrl(ctrl[31]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_32(.inData_0(wireIn[64]), .inData_1(wireIn[65]), .outData_0(wireOut[64]), .outData_1(wireOut[65]), .ctrl(ctrl[32]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_33(.inData_0(wireIn[66]), .inData_1(wireIn[67]), .outData_0(wireOut[66]), .outData_1(wireOut[67]), .ctrl(ctrl[33]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_34(.inData_0(wireIn[68]), .inData_1(wireIn[69]), .outData_0(wireOut[68]), .outData_1(wireOut[69]), .ctrl(ctrl[34]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_35(.inData_0(wireIn[70]), .inData_1(wireIn[71]), .outData_0(wireOut[70]), .outData_1(wireOut[71]), .ctrl(ctrl[35]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_36(.inData_0(wireIn[72]), .inData_1(wireIn[73]), .outData_0(wireOut[72]), .outData_1(wireOut[73]), .ctrl(ctrl[36]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_37(.inData_0(wireIn[74]), .inData_1(wireIn[75]), .outData_0(wireOut[74]), .outData_1(wireOut[75]), .ctrl(ctrl[37]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_38(.inData_0(wireIn[76]), .inData_1(wireIn[77]), .outData_0(wireOut[76]), .outData_1(wireOut[77]), .ctrl(ctrl[38]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_39(.inData_0(wireIn[78]), .inData_1(wireIn[79]), .outData_0(wireOut[78]), .outData_1(wireOut[79]), .ctrl(ctrl[39]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_40(.inData_0(wireIn[80]), .inData_1(wireIn[81]), .outData_0(wireOut[80]), .outData_1(wireOut[81]), .ctrl(ctrl[40]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_41(.inData_0(wireIn[82]), .inData_1(wireIn[83]), .outData_0(wireOut[82]), .outData_1(wireOut[83]), .ctrl(ctrl[41]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_42(.inData_0(wireIn[84]), .inData_1(wireIn[85]), .outData_0(wireOut[84]), .outData_1(wireOut[85]), .ctrl(ctrl[42]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_43(.inData_0(wireIn[86]), .inData_1(wireIn[87]), .outData_0(wireOut[86]), .outData_1(wireOut[87]), .ctrl(ctrl[43]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_44(.inData_0(wireIn[88]), .inData_1(wireIn[89]), .outData_0(wireOut[88]), .outData_1(wireOut[89]), .ctrl(ctrl[44]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_45(.inData_0(wireIn[90]), .inData_1(wireIn[91]), .outData_0(wireOut[90]), .outData_1(wireOut[91]), .ctrl(ctrl[45]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_46(.inData_0(wireIn[92]), .inData_1(wireIn[93]), .outData_0(wireOut[92]), .outData_1(wireOut[93]), .ctrl(ctrl[46]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_47(.inData_0(wireIn[94]), .inData_1(wireIn[95]), .outData_0(wireOut[94]), .outData_1(wireOut[95]), .ctrl(ctrl[47]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_48(.inData_0(wireIn[96]), .inData_1(wireIn[97]), .outData_0(wireOut[96]), .outData_1(wireOut[97]), .ctrl(ctrl[48]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_49(.inData_0(wireIn[98]), .inData_1(wireIn[99]), .outData_0(wireOut[98]), .outData_1(wireOut[99]), .ctrl(ctrl[49]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_50(.inData_0(wireIn[100]), .inData_1(wireIn[101]), .outData_0(wireOut[100]), .outData_1(wireOut[101]), .ctrl(ctrl[50]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_51(.inData_0(wireIn[102]), .inData_1(wireIn[103]), .outData_0(wireOut[102]), .outData_1(wireOut[103]), .ctrl(ctrl[51]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_52(.inData_0(wireIn[104]), .inData_1(wireIn[105]), .outData_0(wireOut[104]), .outData_1(wireOut[105]), .ctrl(ctrl[52]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_53(.inData_0(wireIn[106]), .inData_1(wireIn[107]), .outData_0(wireOut[106]), .outData_1(wireOut[107]), .ctrl(ctrl[53]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_54(.inData_0(wireIn[108]), .inData_1(wireIn[109]), .outData_0(wireOut[108]), .outData_1(wireOut[109]), .ctrl(ctrl[54]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_55(.inData_0(wireIn[110]), .inData_1(wireIn[111]), .outData_0(wireOut[110]), .outData_1(wireOut[111]), .ctrl(ctrl[55]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_56(.inData_0(wireIn[112]), .inData_1(wireIn[113]), .outData_0(wireOut[112]), .outData_1(wireOut[113]), .ctrl(ctrl[56]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_57(.inData_0(wireIn[114]), .inData_1(wireIn[115]), .outData_0(wireOut[114]), .outData_1(wireOut[115]), .ctrl(ctrl[57]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_58(.inData_0(wireIn[116]), .inData_1(wireIn[117]), .outData_0(wireOut[116]), .outData_1(wireOut[117]), .ctrl(ctrl[58]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_59(.inData_0(wireIn[118]), .inData_1(wireIn[119]), .outData_0(wireOut[118]), .outData_1(wireOut[119]), .ctrl(ctrl[59]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_60(.inData_0(wireIn[120]), .inData_1(wireIn[121]), .outData_0(wireOut[120]), .outData_1(wireOut[121]), .ctrl(ctrl[60]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_61(.inData_0(wireIn[122]), .inData_1(wireIn[123]), .outData_0(wireOut[122]), .outData_1(wireOut[123]), .ctrl(ctrl[61]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_62(.inData_0(wireIn[124]), .inData_1(wireIn[125]), .outData_0(wireOut[124]), .outData_1(wireOut[125]), .ctrl(ctrl[62]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_63(.inData_0(wireIn[126]), .inData_1(wireIn[127]), .outData_0(wireOut[126]), .outData_1(wireOut[127]), .ctrl(ctrl[63]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_64(.inData_0(wireIn[128]), .inData_1(wireIn[129]), .outData_0(wireOut[128]), .outData_1(wireOut[129]), .ctrl(ctrl[64]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_65(.inData_0(wireIn[130]), .inData_1(wireIn[131]), .outData_0(wireOut[130]), .outData_1(wireOut[131]), .ctrl(ctrl[65]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_66(.inData_0(wireIn[132]), .inData_1(wireIn[133]), .outData_0(wireOut[132]), .outData_1(wireOut[133]), .ctrl(ctrl[66]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_67(.inData_0(wireIn[134]), .inData_1(wireIn[135]), .outData_0(wireOut[134]), .outData_1(wireOut[135]), .ctrl(ctrl[67]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_68(.inData_0(wireIn[136]), .inData_1(wireIn[137]), .outData_0(wireOut[136]), .outData_1(wireOut[137]), .ctrl(ctrl[68]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_69(.inData_0(wireIn[138]), .inData_1(wireIn[139]), .outData_0(wireOut[138]), .outData_1(wireOut[139]), .ctrl(ctrl[69]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_70(.inData_0(wireIn[140]), .inData_1(wireIn[141]), .outData_0(wireOut[140]), .outData_1(wireOut[141]), .ctrl(ctrl[70]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_71(.inData_0(wireIn[142]), .inData_1(wireIn[143]), .outData_0(wireOut[142]), .outData_1(wireOut[143]), .ctrl(ctrl[71]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_72(.inData_0(wireIn[144]), .inData_1(wireIn[145]), .outData_0(wireOut[144]), .outData_1(wireOut[145]), .ctrl(ctrl[72]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_73(.inData_0(wireIn[146]), .inData_1(wireIn[147]), .outData_0(wireOut[146]), .outData_1(wireOut[147]), .ctrl(ctrl[73]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_74(.inData_0(wireIn[148]), .inData_1(wireIn[149]), .outData_0(wireOut[148]), .outData_1(wireOut[149]), .ctrl(ctrl[74]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_75(.inData_0(wireIn[150]), .inData_1(wireIn[151]), .outData_0(wireOut[150]), .outData_1(wireOut[151]), .ctrl(ctrl[75]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_76(.inData_0(wireIn[152]), .inData_1(wireIn[153]), .outData_0(wireOut[152]), .outData_1(wireOut[153]), .ctrl(ctrl[76]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_77(.inData_0(wireIn[154]), .inData_1(wireIn[155]), .outData_0(wireOut[154]), .outData_1(wireOut[155]), .ctrl(ctrl[77]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_78(.inData_0(wireIn[156]), .inData_1(wireIn[157]), .outData_0(wireOut[156]), .outData_1(wireOut[157]), .ctrl(ctrl[78]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_79(.inData_0(wireIn[158]), .inData_1(wireIn[159]), .outData_0(wireOut[158]), .outData_1(wireOut[159]), .ctrl(ctrl[79]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_80(.inData_0(wireIn[160]), .inData_1(wireIn[161]), .outData_0(wireOut[160]), .outData_1(wireOut[161]), .ctrl(ctrl[80]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_81(.inData_0(wireIn[162]), .inData_1(wireIn[163]), .outData_0(wireOut[162]), .outData_1(wireOut[163]), .ctrl(ctrl[81]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_82(.inData_0(wireIn[164]), .inData_1(wireIn[165]), .outData_0(wireOut[164]), .outData_1(wireOut[165]), .ctrl(ctrl[82]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_83(.inData_0(wireIn[166]), .inData_1(wireIn[167]), .outData_0(wireOut[166]), .outData_1(wireOut[167]), .ctrl(ctrl[83]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_84(.inData_0(wireIn[168]), .inData_1(wireIn[169]), .outData_0(wireOut[168]), .outData_1(wireOut[169]), .ctrl(ctrl[84]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_85(.inData_0(wireIn[170]), .inData_1(wireIn[171]), .outData_0(wireOut[170]), .outData_1(wireOut[171]), .ctrl(ctrl[85]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_86(.inData_0(wireIn[172]), .inData_1(wireIn[173]), .outData_0(wireOut[172]), .outData_1(wireOut[173]), .ctrl(ctrl[86]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_87(.inData_0(wireIn[174]), .inData_1(wireIn[175]), .outData_0(wireOut[174]), .outData_1(wireOut[175]), .ctrl(ctrl[87]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_88(.inData_0(wireIn[176]), .inData_1(wireIn[177]), .outData_0(wireOut[176]), .outData_1(wireOut[177]), .ctrl(ctrl[88]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_89(.inData_0(wireIn[178]), .inData_1(wireIn[179]), .outData_0(wireOut[178]), .outData_1(wireOut[179]), .ctrl(ctrl[89]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_90(.inData_0(wireIn[180]), .inData_1(wireIn[181]), .outData_0(wireOut[180]), .outData_1(wireOut[181]), .ctrl(ctrl[90]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_91(.inData_0(wireIn[182]), .inData_1(wireIn[183]), .outData_0(wireOut[182]), .outData_1(wireOut[183]), .ctrl(ctrl[91]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_92(.inData_0(wireIn[184]), .inData_1(wireIn[185]), .outData_0(wireOut[184]), .outData_1(wireOut[185]), .ctrl(ctrl[92]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_93(.inData_0(wireIn[186]), .inData_1(wireIn[187]), .outData_0(wireOut[186]), .outData_1(wireOut[187]), .ctrl(ctrl[93]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_94(.inData_0(wireIn[188]), .inData_1(wireIn[189]), .outData_0(wireOut[188]), .outData_1(wireOut[189]), .ctrl(ctrl[94]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_95(.inData_0(wireIn[190]), .inData_1(wireIn[191]), .outData_0(wireOut[190]), .outData_1(wireOut[191]), .ctrl(ctrl[95]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_96(.inData_0(wireIn[192]), .inData_1(wireIn[193]), .outData_0(wireOut[192]), .outData_1(wireOut[193]), .ctrl(ctrl[96]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_97(.inData_0(wireIn[194]), .inData_1(wireIn[195]), .outData_0(wireOut[194]), .outData_1(wireOut[195]), .ctrl(ctrl[97]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_98(.inData_0(wireIn[196]), .inData_1(wireIn[197]), .outData_0(wireOut[196]), .outData_1(wireOut[197]), .ctrl(ctrl[98]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_99(.inData_0(wireIn[198]), .inData_1(wireIn[199]), .outData_0(wireOut[198]), .outData_1(wireOut[199]), .ctrl(ctrl[99]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_100(.inData_0(wireIn[200]), .inData_1(wireIn[201]), .outData_0(wireOut[200]), .outData_1(wireOut[201]), .ctrl(ctrl[100]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_101(.inData_0(wireIn[202]), .inData_1(wireIn[203]), .outData_0(wireOut[202]), .outData_1(wireOut[203]), .ctrl(ctrl[101]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_102(.inData_0(wireIn[204]), .inData_1(wireIn[205]), .outData_0(wireOut[204]), .outData_1(wireOut[205]), .ctrl(ctrl[102]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_103(.inData_0(wireIn[206]), .inData_1(wireIn[207]), .outData_0(wireOut[206]), .outData_1(wireOut[207]), .ctrl(ctrl[103]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_104(.inData_0(wireIn[208]), .inData_1(wireIn[209]), .outData_0(wireOut[208]), .outData_1(wireOut[209]), .ctrl(ctrl[104]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_105(.inData_0(wireIn[210]), .inData_1(wireIn[211]), .outData_0(wireOut[210]), .outData_1(wireOut[211]), .ctrl(ctrl[105]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_106(.inData_0(wireIn[212]), .inData_1(wireIn[213]), .outData_0(wireOut[212]), .outData_1(wireOut[213]), .ctrl(ctrl[106]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_107(.inData_0(wireIn[214]), .inData_1(wireIn[215]), .outData_0(wireOut[214]), .outData_1(wireOut[215]), .ctrl(ctrl[107]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_108(.inData_0(wireIn[216]), .inData_1(wireIn[217]), .outData_0(wireOut[216]), .outData_1(wireOut[217]), .ctrl(ctrl[108]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_109(.inData_0(wireIn[218]), .inData_1(wireIn[219]), .outData_0(wireOut[218]), .outData_1(wireOut[219]), .ctrl(ctrl[109]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_110(.inData_0(wireIn[220]), .inData_1(wireIn[221]), .outData_0(wireOut[220]), .outData_1(wireOut[221]), .ctrl(ctrl[110]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_111(.inData_0(wireIn[222]), .inData_1(wireIn[223]), .outData_0(wireOut[222]), .outData_1(wireOut[223]), .ctrl(ctrl[111]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_112(.inData_0(wireIn[224]), .inData_1(wireIn[225]), .outData_0(wireOut[224]), .outData_1(wireOut[225]), .ctrl(ctrl[112]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_113(.inData_0(wireIn[226]), .inData_1(wireIn[227]), .outData_0(wireOut[226]), .outData_1(wireOut[227]), .ctrl(ctrl[113]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_114(.inData_0(wireIn[228]), .inData_1(wireIn[229]), .outData_0(wireOut[228]), .outData_1(wireOut[229]), .ctrl(ctrl[114]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_115(.inData_0(wireIn[230]), .inData_1(wireIn[231]), .outData_0(wireOut[230]), .outData_1(wireOut[231]), .ctrl(ctrl[115]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_116(.inData_0(wireIn[232]), .inData_1(wireIn[233]), .outData_0(wireOut[232]), .outData_1(wireOut[233]), .ctrl(ctrl[116]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_117(.inData_0(wireIn[234]), .inData_1(wireIn[235]), .outData_0(wireOut[234]), .outData_1(wireOut[235]), .ctrl(ctrl[117]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_118(.inData_0(wireIn[236]), .inData_1(wireIn[237]), .outData_0(wireOut[236]), .outData_1(wireOut[237]), .ctrl(ctrl[118]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_119(.inData_0(wireIn[238]), .inData_1(wireIn[239]), .outData_0(wireOut[238]), .outData_1(wireOut[239]), .ctrl(ctrl[119]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_120(.inData_0(wireIn[240]), .inData_1(wireIn[241]), .outData_0(wireOut[240]), .outData_1(wireOut[241]), .ctrl(ctrl[120]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_121(.inData_0(wireIn[242]), .inData_1(wireIn[243]), .outData_0(wireOut[242]), .outData_1(wireOut[243]), .ctrl(ctrl[121]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_122(.inData_0(wireIn[244]), .inData_1(wireIn[245]), .outData_0(wireOut[244]), .outData_1(wireOut[245]), .ctrl(ctrl[122]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_123(.inData_0(wireIn[246]), .inData_1(wireIn[247]), .outData_0(wireOut[246]), .outData_1(wireOut[247]), .ctrl(ctrl[123]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_124(.inData_0(wireIn[248]), .inData_1(wireIn[249]), .outData_0(wireOut[248]), .outData_1(wireOut[249]), .ctrl(ctrl[124]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_125(.inData_0(wireIn[250]), .inData_1(wireIn[251]), .outData_0(wireOut[250]), .outData_1(wireOut[251]), .ctrl(ctrl[125]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_126(.inData_0(wireIn[252]), .inData_1(wireIn[253]), .outData_0(wireOut[252]), .outData_1(wireOut[253]), .ctrl(ctrl[126]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_127(.inData_0(wireIn[254]), .inData_1(wireIn[255]), .outData_0(wireOut[254]), .outData_1(wireOut[255]), .ctrl(ctrl[127]), .clk(clk), .rst(rst));
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module wireCon_dp256_st0_L(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  assign wireOut[0] = wireIn[0];    
  assign wireOut[1] = wireIn[2];    
  assign wireOut[2] = wireIn[4];    
  assign wireOut[3] = wireIn[6];    
  assign wireOut[4] = wireIn[8];    
  assign wireOut[5] = wireIn[10];    
  assign wireOut[6] = wireIn[12];    
  assign wireOut[7] = wireIn[14];    
  assign wireOut[8] = wireIn[16];    
  assign wireOut[9] = wireIn[18];    
  assign wireOut[10] = wireIn[20];    
  assign wireOut[11] = wireIn[22];    
  assign wireOut[12] = wireIn[24];    
  assign wireOut[13] = wireIn[26];    
  assign wireOut[14] = wireIn[28];    
  assign wireOut[15] = wireIn[30];    
  assign wireOut[16] = wireIn[32];    
  assign wireOut[17] = wireIn[34];    
  assign wireOut[18] = wireIn[36];    
  assign wireOut[19] = wireIn[38];    
  assign wireOut[20] = wireIn[40];    
  assign wireOut[21] = wireIn[42];    
  assign wireOut[22] = wireIn[44];    
  assign wireOut[23] = wireIn[46];    
  assign wireOut[24] = wireIn[48];    
  assign wireOut[25] = wireIn[50];    
  assign wireOut[26] = wireIn[52];    
  assign wireOut[27] = wireIn[54];    
  assign wireOut[28] = wireIn[56];    
  assign wireOut[29] = wireIn[58];    
  assign wireOut[30] = wireIn[60];    
  assign wireOut[31] = wireIn[62];    
  assign wireOut[32] = wireIn[64];    
  assign wireOut[33] = wireIn[66];    
  assign wireOut[34] = wireIn[68];    
  assign wireOut[35] = wireIn[70];    
  assign wireOut[36] = wireIn[72];    
  assign wireOut[37] = wireIn[74];    
  assign wireOut[38] = wireIn[76];    
  assign wireOut[39] = wireIn[78];    
  assign wireOut[40] = wireIn[80];    
  assign wireOut[41] = wireIn[82];    
  assign wireOut[42] = wireIn[84];    
  assign wireOut[43] = wireIn[86];    
  assign wireOut[44] = wireIn[88];    
  assign wireOut[45] = wireIn[90];    
  assign wireOut[46] = wireIn[92];    
  assign wireOut[47] = wireIn[94];    
  assign wireOut[48] = wireIn[96];    
  assign wireOut[49] = wireIn[98];    
  assign wireOut[50] = wireIn[100];    
  assign wireOut[51] = wireIn[102];    
  assign wireOut[52] = wireIn[104];    
  assign wireOut[53] = wireIn[106];    
  assign wireOut[54] = wireIn[108];    
  assign wireOut[55] = wireIn[110];    
  assign wireOut[56] = wireIn[112];    
  assign wireOut[57] = wireIn[114];    
  assign wireOut[58] = wireIn[116];    
  assign wireOut[59] = wireIn[118];    
  assign wireOut[60] = wireIn[120];    
  assign wireOut[61] = wireIn[122];    
  assign wireOut[62] = wireIn[124];    
  assign wireOut[63] = wireIn[126];    
  assign wireOut[64] = wireIn[128];    
  assign wireOut[65] = wireIn[130];    
  assign wireOut[66] = wireIn[132];    
  assign wireOut[67] = wireIn[134];    
  assign wireOut[68] = wireIn[136];    
  assign wireOut[69] = wireIn[138];    
  assign wireOut[70] = wireIn[140];    
  assign wireOut[71] = wireIn[142];    
  assign wireOut[72] = wireIn[144];    
  assign wireOut[73] = wireIn[146];    
  assign wireOut[74] = wireIn[148];    
  assign wireOut[75] = wireIn[150];    
  assign wireOut[76] = wireIn[152];    
  assign wireOut[77] = wireIn[154];    
  assign wireOut[78] = wireIn[156];    
  assign wireOut[79] = wireIn[158];    
  assign wireOut[80] = wireIn[160];    
  assign wireOut[81] = wireIn[162];    
  assign wireOut[82] = wireIn[164];    
  assign wireOut[83] = wireIn[166];    
  assign wireOut[84] = wireIn[168];    
  assign wireOut[85] = wireIn[170];    
  assign wireOut[86] = wireIn[172];    
  assign wireOut[87] = wireIn[174];    
  assign wireOut[88] = wireIn[176];    
  assign wireOut[89] = wireIn[178];    
  assign wireOut[90] = wireIn[180];    
  assign wireOut[91] = wireIn[182];    
  assign wireOut[92] = wireIn[184];    
  assign wireOut[93] = wireIn[186];    
  assign wireOut[94] = wireIn[188];    
  assign wireOut[95] = wireIn[190];    
  assign wireOut[96] = wireIn[192];    
  assign wireOut[97] = wireIn[194];    
  assign wireOut[98] = wireIn[196];    
  assign wireOut[99] = wireIn[198];    
  assign wireOut[100] = wireIn[200];    
  assign wireOut[101] = wireIn[202];    
  assign wireOut[102] = wireIn[204];    
  assign wireOut[103] = wireIn[206];    
  assign wireOut[104] = wireIn[208];    
  assign wireOut[105] = wireIn[210];    
  assign wireOut[106] = wireIn[212];    
  assign wireOut[107] = wireIn[214];    
  assign wireOut[108] = wireIn[216];    
  assign wireOut[109] = wireIn[218];    
  assign wireOut[110] = wireIn[220];    
  assign wireOut[111] = wireIn[222];    
  assign wireOut[112] = wireIn[224];    
  assign wireOut[113] = wireIn[226];    
  assign wireOut[114] = wireIn[228];    
  assign wireOut[115] = wireIn[230];    
  assign wireOut[116] = wireIn[232];    
  assign wireOut[117] = wireIn[234];    
  assign wireOut[118] = wireIn[236];    
  assign wireOut[119] = wireIn[238];    
  assign wireOut[120] = wireIn[240];    
  assign wireOut[121] = wireIn[242];    
  assign wireOut[122] = wireIn[244];    
  assign wireOut[123] = wireIn[246];    
  assign wireOut[124] = wireIn[248];    
  assign wireOut[125] = wireIn[250];    
  assign wireOut[126] = wireIn[252];    
  assign wireOut[127] = wireIn[254];    
  assign wireOut[128] = wireIn[1];    
  assign wireOut[129] = wireIn[3];    
  assign wireOut[130] = wireIn[5];    
  assign wireOut[131] = wireIn[7];    
  assign wireOut[132] = wireIn[9];    
  assign wireOut[133] = wireIn[11];    
  assign wireOut[134] = wireIn[13];    
  assign wireOut[135] = wireIn[15];    
  assign wireOut[136] = wireIn[17];    
  assign wireOut[137] = wireIn[19];    
  assign wireOut[138] = wireIn[21];    
  assign wireOut[139] = wireIn[23];    
  assign wireOut[140] = wireIn[25];    
  assign wireOut[141] = wireIn[27];    
  assign wireOut[142] = wireIn[29];    
  assign wireOut[143] = wireIn[31];    
  assign wireOut[144] = wireIn[33];    
  assign wireOut[145] = wireIn[35];    
  assign wireOut[146] = wireIn[37];    
  assign wireOut[147] = wireIn[39];    
  assign wireOut[148] = wireIn[41];    
  assign wireOut[149] = wireIn[43];    
  assign wireOut[150] = wireIn[45];    
  assign wireOut[151] = wireIn[47];    
  assign wireOut[152] = wireIn[49];    
  assign wireOut[153] = wireIn[51];    
  assign wireOut[154] = wireIn[53];    
  assign wireOut[155] = wireIn[55];    
  assign wireOut[156] = wireIn[57];    
  assign wireOut[157] = wireIn[59];    
  assign wireOut[158] = wireIn[61];    
  assign wireOut[159] = wireIn[63];    
  assign wireOut[160] = wireIn[65];    
  assign wireOut[161] = wireIn[67];    
  assign wireOut[162] = wireIn[69];    
  assign wireOut[163] = wireIn[71];    
  assign wireOut[164] = wireIn[73];    
  assign wireOut[165] = wireIn[75];    
  assign wireOut[166] = wireIn[77];    
  assign wireOut[167] = wireIn[79];    
  assign wireOut[168] = wireIn[81];    
  assign wireOut[169] = wireIn[83];    
  assign wireOut[170] = wireIn[85];    
  assign wireOut[171] = wireIn[87];    
  assign wireOut[172] = wireIn[89];    
  assign wireOut[173] = wireIn[91];    
  assign wireOut[174] = wireIn[93];    
  assign wireOut[175] = wireIn[95];    
  assign wireOut[176] = wireIn[97];    
  assign wireOut[177] = wireIn[99];    
  assign wireOut[178] = wireIn[101];    
  assign wireOut[179] = wireIn[103];    
  assign wireOut[180] = wireIn[105];    
  assign wireOut[181] = wireIn[107];    
  assign wireOut[182] = wireIn[109];    
  assign wireOut[183] = wireIn[111];    
  assign wireOut[184] = wireIn[113];    
  assign wireOut[185] = wireIn[115];    
  assign wireOut[186] = wireIn[117];    
  assign wireOut[187] = wireIn[119];    
  assign wireOut[188] = wireIn[121];    
  assign wireOut[189] = wireIn[123];    
  assign wireOut[190] = wireIn[125];    
  assign wireOut[191] = wireIn[127];    
  assign wireOut[192] = wireIn[129];    
  assign wireOut[193] = wireIn[131];    
  assign wireOut[194] = wireIn[133];    
  assign wireOut[195] = wireIn[135];    
  assign wireOut[196] = wireIn[137];    
  assign wireOut[197] = wireIn[139];    
  assign wireOut[198] = wireIn[141];    
  assign wireOut[199] = wireIn[143];    
  assign wireOut[200] = wireIn[145];    
  assign wireOut[201] = wireIn[147];    
  assign wireOut[202] = wireIn[149];    
  assign wireOut[203] = wireIn[151];    
  assign wireOut[204] = wireIn[153];    
  assign wireOut[205] = wireIn[155];    
  assign wireOut[206] = wireIn[157];    
  assign wireOut[207] = wireIn[159];    
  assign wireOut[208] = wireIn[161];    
  assign wireOut[209] = wireIn[163];    
  assign wireOut[210] = wireIn[165];    
  assign wireOut[211] = wireIn[167];    
  assign wireOut[212] = wireIn[169];    
  assign wireOut[213] = wireIn[171];    
  assign wireOut[214] = wireIn[173];    
  assign wireOut[215] = wireIn[175];    
  assign wireOut[216] = wireIn[177];    
  assign wireOut[217] = wireIn[179];    
  assign wireOut[218] = wireIn[181];    
  assign wireOut[219] = wireIn[183];    
  assign wireOut[220] = wireIn[185];    
  assign wireOut[221] = wireIn[187];    
  assign wireOut[222] = wireIn[189];    
  assign wireOut[223] = wireIn[191];    
  assign wireOut[224] = wireIn[193];    
  assign wireOut[225] = wireIn[195];    
  assign wireOut[226] = wireIn[197];    
  assign wireOut[227] = wireIn[199];    
  assign wireOut[228] = wireIn[201];    
  assign wireOut[229] = wireIn[203];    
  assign wireOut[230] = wireIn[205];    
  assign wireOut[231] = wireIn[207];    
  assign wireOut[232] = wireIn[209];    
  assign wireOut[233] = wireIn[211];    
  assign wireOut[234] = wireIn[213];    
  assign wireOut[235] = wireIn[215];    
  assign wireOut[236] = wireIn[217];    
  assign wireOut[237] = wireIn[219];    
  assign wireOut[238] = wireIn[221];    
  assign wireOut[239] = wireIn[223];    
  assign wireOut[240] = wireIn[225];    
  assign wireOut[241] = wireIn[227];    
  assign wireOut[242] = wireIn[229];    
  assign wireOut[243] = wireIn[231];    
  assign wireOut[244] = wireIn[233];    
  assign wireOut[245] = wireIn[235];    
  assign wireOut[246] = wireIn[237];    
  assign wireOut[247] = wireIn[239];    
  assign wireOut[248] = wireIn[241];    
  assign wireOut[249] = wireIn[243];    
  assign wireOut[250] = wireIn[245];    
  assign wireOut[251] = wireIn[247];    
  assign wireOut[252] = wireIn[249];    
  assign wireOut[253] = wireIn[251];    
  assign wireOut[254] = wireIn[253];    
  assign wireOut[255] = wireIn[255];    
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module switches_stage_st1_0_L(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
ctrl,                            
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;                   
  input [128-1:0] ctrl;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  switch_2_2 switch_inst_0(.inData_0(wireIn[0]), .inData_1(wireIn[1]), .outData_0(wireOut[0]), .outData_1(wireOut[1]), .ctrl(ctrl[0]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_1(.inData_0(wireIn[2]), .inData_1(wireIn[3]), .outData_0(wireOut[2]), .outData_1(wireOut[3]), .ctrl(ctrl[1]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_2(.inData_0(wireIn[4]), .inData_1(wireIn[5]), .outData_0(wireOut[4]), .outData_1(wireOut[5]), .ctrl(ctrl[2]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_3(.inData_0(wireIn[6]), .inData_1(wireIn[7]), .outData_0(wireOut[6]), .outData_1(wireOut[7]), .ctrl(ctrl[3]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_4(.inData_0(wireIn[8]), .inData_1(wireIn[9]), .outData_0(wireOut[8]), .outData_1(wireOut[9]), .ctrl(ctrl[4]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_5(.inData_0(wireIn[10]), .inData_1(wireIn[11]), .outData_0(wireOut[10]), .outData_1(wireOut[11]), .ctrl(ctrl[5]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_6(.inData_0(wireIn[12]), .inData_1(wireIn[13]), .outData_0(wireOut[12]), .outData_1(wireOut[13]), .ctrl(ctrl[6]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_7(.inData_0(wireIn[14]), .inData_1(wireIn[15]), .outData_0(wireOut[14]), .outData_1(wireOut[15]), .ctrl(ctrl[7]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_8(.inData_0(wireIn[16]), .inData_1(wireIn[17]), .outData_0(wireOut[16]), .outData_1(wireOut[17]), .ctrl(ctrl[8]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_9(.inData_0(wireIn[18]), .inData_1(wireIn[19]), .outData_0(wireOut[18]), .outData_1(wireOut[19]), .ctrl(ctrl[9]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_10(.inData_0(wireIn[20]), .inData_1(wireIn[21]), .outData_0(wireOut[20]), .outData_1(wireOut[21]), .ctrl(ctrl[10]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_11(.inData_0(wireIn[22]), .inData_1(wireIn[23]), .outData_0(wireOut[22]), .outData_1(wireOut[23]), .ctrl(ctrl[11]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_12(.inData_0(wireIn[24]), .inData_1(wireIn[25]), .outData_0(wireOut[24]), .outData_1(wireOut[25]), .ctrl(ctrl[12]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_13(.inData_0(wireIn[26]), .inData_1(wireIn[27]), .outData_0(wireOut[26]), .outData_1(wireOut[27]), .ctrl(ctrl[13]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_14(.inData_0(wireIn[28]), .inData_1(wireIn[29]), .outData_0(wireOut[28]), .outData_1(wireOut[29]), .ctrl(ctrl[14]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_15(.inData_0(wireIn[30]), .inData_1(wireIn[31]), .outData_0(wireOut[30]), .outData_1(wireOut[31]), .ctrl(ctrl[15]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_16(.inData_0(wireIn[32]), .inData_1(wireIn[33]), .outData_0(wireOut[32]), .outData_1(wireOut[33]), .ctrl(ctrl[16]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_17(.inData_0(wireIn[34]), .inData_1(wireIn[35]), .outData_0(wireOut[34]), .outData_1(wireOut[35]), .ctrl(ctrl[17]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_18(.inData_0(wireIn[36]), .inData_1(wireIn[37]), .outData_0(wireOut[36]), .outData_1(wireOut[37]), .ctrl(ctrl[18]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_19(.inData_0(wireIn[38]), .inData_1(wireIn[39]), .outData_0(wireOut[38]), .outData_1(wireOut[39]), .ctrl(ctrl[19]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_20(.inData_0(wireIn[40]), .inData_1(wireIn[41]), .outData_0(wireOut[40]), .outData_1(wireOut[41]), .ctrl(ctrl[20]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_21(.inData_0(wireIn[42]), .inData_1(wireIn[43]), .outData_0(wireOut[42]), .outData_1(wireOut[43]), .ctrl(ctrl[21]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_22(.inData_0(wireIn[44]), .inData_1(wireIn[45]), .outData_0(wireOut[44]), .outData_1(wireOut[45]), .ctrl(ctrl[22]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_23(.inData_0(wireIn[46]), .inData_1(wireIn[47]), .outData_0(wireOut[46]), .outData_1(wireOut[47]), .ctrl(ctrl[23]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_24(.inData_0(wireIn[48]), .inData_1(wireIn[49]), .outData_0(wireOut[48]), .outData_1(wireOut[49]), .ctrl(ctrl[24]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_25(.inData_0(wireIn[50]), .inData_1(wireIn[51]), .outData_0(wireOut[50]), .outData_1(wireOut[51]), .ctrl(ctrl[25]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_26(.inData_0(wireIn[52]), .inData_1(wireIn[53]), .outData_0(wireOut[52]), .outData_1(wireOut[53]), .ctrl(ctrl[26]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_27(.inData_0(wireIn[54]), .inData_1(wireIn[55]), .outData_0(wireOut[54]), .outData_1(wireOut[55]), .ctrl(ctrl[27]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_28(.inData_0(wireIn[56]), .inData_1(wireIn[57]), .outData_0(wireOut[56]), .outData_1(wireOut[57]), .ctrl(ctrl[28]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_29(.inData_0(wireIn[58]), .inData_1(wireIn[59]), .outData_0(wireOut[58]), .outData_1(wireOut[59]), .ctrl(ctrl[29]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_30(.inData_0(wireIn[60]), .inData_1(wireIn[61]), .outData_0(wireOut[60]), .outData_1(wireOut[61]), .ctrl(ctrl[30]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_31(.inData_0(wireIn[62]), .inData_1(wireIn[63]), .outData_0(wireOut[62]), .outData_1(wireOut[63]), .ctrl(ctrl[31]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_32(.inData_0(wireIn[64]), .inData_1(wireIn[65]), .outData_0(wireOut[64]), .outData_1(wireOut[65]), .ctrl(ctrl[32]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_33(.inData_0(wireIn[66]), .inData_1(wireIn[67]), .outData_0(wireOut[66]), .outData_1(wireOut[67]), .ctrl(ctrl[33]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_34(.inData_0(wireIn[68]), .inData_1(wireIn[69]), .outData_0(wireOut[68]), .outData_1(wireOut[69]), .ctrl(ctrl[34]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_35(.inData_0(wireIn[70]), .inData_1(wireIn[71]), .outData_0(wireOut[70]), .outData_1(wireOut[71]), .ctrl(ctrl[35]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_36(.inData_0(wireIn[72]), .inData_1(wireIn[73]), .outData_0(wireOut[72]), .outData_1(wireOut[73]), .ctrl(ctrl[36]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_37(.inData_0(wireIn[74]), .inData_1(wireIn[75]), .outData_0(wireOut[74]), .outData_1(wireOut[75]), .ctrl(ctrl[37]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_38(.inData_0(wireIn[76]), .inData_1(wireIn[77]), .outData_0(wireOut[76]), .outData_1(wireOut[77]), .ctrl(ctrl[38]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_39(.inData_0(wireIn[78]), .inData_1(wireIn[79]), .outData_0(wireOut[78]), .outData_1(wireOut[79]), .ctrl(ctrl[39]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_40(.inData_0(wireIn[80]), .inData_1(wireIn[81]), .outData_0(wireOut[80]), .outData_1(wireOut[81]), .ctrl(ctrl[40]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_41(.inData_0(wireIn[82]), .inData_1(wireIn[83]), .outData_0(wireOut[82]), .outData_1(wireOut[83]), .ctrl(ctrl[41]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_42(.inData_0(wireIn[84]), .inData_1(wireIn[85]), .outData_0(wireOut[84]), .outData_1(wireOut[85]), .ctrl(ctrl[42]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_43(.inData_0(wireIn[86]), .inData_1(wireIn[87]), .outData_0(wireOut[86]), .outData_1(wireOut[87]), .ctrl(ctrl[43]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_44(.inData_0(wireIn[88]), .inData_1(wireIn[89]), .outData_0(wireOut[88]), .outData_1(wireOut[89]), .ctrl(ctrl[44]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_45(.inData_0(wireIn[90]), .inData_1(wireIn[91]), .outData_0(wireOut[90]), .outData_1(wireOut[91]), .ctrl(ctrl[45]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_46(.inData_0(wireIn[92]), .inData_1(wireIn[93]), .outData_0(wireOut[92]), .outData_1(wireOut[93]), .ctrl(ctrl[46]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_47(.inData_0(wireIn[94]), .inData_1(wireIn[95]), .outData_0(wireOut[94]), .outData_1(wireOut[95]), .ctrl(ctrl[47]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_48(.inData_0(wireIn[96]), .inData_1(wireIn[97]), .outData_0(wireOut[96]), .outData_1(wireOut[97]), .ctrl(ctrl[48]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_49(.inData_0(wireIn[98]), .inData_1(wireIn[99]), .outData_0(wireOut[98]), .outData_1(wireOut[99]), .ctrl(ctrl[49]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_50(.inData_0(wireIn[100]), .inData_1(wireIn[101]), .outData_0(wireOut[100]), .outData_1(wireOut[101]), .ctrl(ctrl[50]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_51(.inData_0(wireIn[102]), .inData_1(wireIn[103]), .outData_0(wireOut[102]), .outData_1(wireOut[103]), .ctrl(ctrl[51]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_52(.inData_0(wireIn[104]), .inData_1(wireIn[105]), .outData_0(wireOut[104]), .outData_1(wireOut[105]), .ctrl(ctrl[52]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_53(.inData_0(wireIn[106]), .inData_1(wireIn[107]), .outData_0(wireOut[106]), .outData_1(wireOut[107]), .ctrl(ctrl[53]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_54(.inData_0(wireIn[108]), .inData_1(wireIn[109]), .outData_0(wireOut[108]), .outData_1(wireOut[109]), .ctrl(ctrl[54]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_55(.inData_0(wireIn[110]), .inData_1(wireIn[111]), .outData_0(wireOut[110]), .outData_1(wireOut[111]), .ctrl(ctrl[55]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_56(.inData_0(wireIn[112]), .inData_1(wireIn[113]), .outData_0(wireOut[112]), .outData_1(wireOut[113]), .ctrl(ctrl[56]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_57(.inData_0(wireIn[114]), .inData_1(wireIn[115]), .outData_0(wireOut[114]), .outData_1(wireOut[115]), .ctrl(ctrl[57]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_58(.inData_0(wireIn[116]), .inData_1(wireIn[117]), .outData_0(wireOut[116]), .outData_1(wireOut[117]), .ctrl(ctrl[58]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_59(.inData_0(wireIn[118]), .inData_1(wireIn[119]), .outData_0(wireOut[118]), .outData_1(wireOut[119]), .ctrl(ctrl[59]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_60(.inData_0(wireIn[120]), .inData_1(wireIn[121]), .outData_0(wireOut[120]), .outData_1(wireOut[121]), .ctrl(ctrl[60]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_61(.inData_0(wireIn[122]), .inData_1(wireIn[123]), .outData_0(wireOut[122]), .outData_1(wireOut[123]), .ctrl(ctrl[61]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_62(.inData_0(wireIn[124]), .inData_1(wireIn[125]), .outData_0(wireOut[124]), .outData_1(wireOut[125]), .ctrl(ctrl[62]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_63(.inData_0(wireIn[126]), .inData_1(wireIn[127]), .outData_0(wireOut[126]), .outData_1(wireOut[127]), .ctrl(ctrl[63]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_64(.inData_0(wireIn[128]), .inData_1(wireIn[129]), .outData_0(wireOut[128]), .outData_1(wireOut[129]), .ctrl(ctrl[64]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_65(.inData_0(wireIn[130]), .inData_1(wireIn[131]), .outData_0(wireOut[130]), .outData_1(wireOut[131]), .ctrl(ctrl[65]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_66(.inData_0(wireIn[132]), .inData_1(wireIn[133]), .outData_0(wireOut[132]), .outData_1(wireOut[133]), .ctrl(ctrl[66]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_67(.inData_0(wireIn[134]), .inData_1(wireIn[135]), .outData_0(wireOut[134]), .outData_1(wireOut[135]), .ctrl(ctrl[67]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_68(.inData_0(wireIn[136]), .inData_1(wireIn[137]), .outData_0(wireOut[136]), .outData_1(wireOut[137]), .ctrl(ctrl[68]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_69(.inData_0(wireIn[138]), .inData_1(wireIn[139]), .outData_0(wireOut[138]), .outData_1(wireOut[139]), .ctrl(ctrl[69]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_70(.inData_0(wireIn[140]), .inData_1(wireIn[141]), .outData_0(wireOut[140]), .outData_1(wireOut[141]), .ctrl(ctrl[70]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_71(.inData_0(wireIn[142]), .inData_1(wireIn[143]), .outData_0(wireOut[142]), .outData_1(wireOut[143]), .ctrl(ctrl[71]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_72(.inData_0(wireIn[144]), .inData_1(wireIn[145]), .outData_0(wireOut[144]), .outData_1(wireOut[145]), .ctrl(ctrl[72]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_73(.inData_0(wireIn[146]), .inData_1(wireIn[147]), .outData_0(wireOut[146]), .outData_1(wireOut[147]), .ctrl(ctrl[73]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_74(.inData_0(wireIn[148]), .inData_1(wireIn[149]), .outData_0(wireOut[148]), .outData_1(wireOut[149]), .ctrl(ctrl[74]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_75(.inData_0(wireIn[150]), .inData_1(wireIn[151]), .outData_0(wireOut[150]), .outData_1(wireOut[151]), .ctrl(ctrl[75]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_76(.inData_0(wireIn[152]), .inData_1(wireIn[153]), .outData_0(wireOut[152]), .outData_1(wireOut[153]), .ctrl(ctrl[76]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_77(.inData_0(wireIn[154]), .inData_1(wireIn[155]), .outData_0(wireOut[154]), .outData_1(wireOut[155]), .ctrl(ctrl[77]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_78(.inData_0(wireIn[156]), .inData_1(wireIn[157]), .outData_0(wireOut[156]), .outData_1(wireOut[157]), .ctrl(ctrl[78]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_79(.inData_0(wireIn[158]), .inData_1(wireIn[159]), .outData_0(wireOut[158]), .outData_1(wireOut[159]), .ctrl(ctrl[79]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_80(.inData_0(wireIn[160]), .inData_1(wireIn[161]), .outData_0(wireOut[160]), .outData_1(wireOut[161]), .ctrl(ctrl[80]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_81(.inData_0(wireIn[162]), .inData_1(wireIn[163]), .outData_0(wireOut[162]), .outData_1(wireOut[163]), .ctrl(ctrl[81]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_82(.inData_0(wireIn[164]), .inData_1(wireIn[165]), .outData_0(wireOut[164]), .outData_1(wireOut[165]), .ctrl(ctrl[82]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_83(.inData_0(wireIn[166]), .inData_1(wireIn[167]), .outData_0(wireOut[166]), .outData_1(wireOut[167]), .ctrl(ctrl[83]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_84(.inData_0(wireIn[168]), .inData_1(wireIn[169]), .outData_0(wireOut[168]), .outData_1(wireOut[169]), .ctrl(ctrl[84]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_85(.inData_0(wireIn[170]), .inData_1(wireIn[171]), .outData_0(wireOut[170]), .outData_1(wireOut[171]), .ctrl(ctrl[85]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_86(.inData_0(wireIn[172]), .inData_1(wireIn[173]), .outData_0(wireOut[172]), .outData_1(wireOut[173]), .ctrl(ctrl[86]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_87(.inData_0(wireIn[174]), .inData_1(wireIn[175]), .outData_0(wireOut[174]), .outData_1(wireOut[175]), .ctrl(ctrl[87]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_88(.inData_0(wireIn[176]), .inData_1(wireIn[177]), .outData_0(wireOut[176]), .outData_1(wireOut[177]), .ctrl(ctrl[88]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_89(.inData_0(wireIn[178]), .inData_1(wireIn[179]), .outData_0(wireOut[178]), .outData_1(wireOut[179]), .ctrl(ctrl[89]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_90(.inData_0(wireIn[180]), .inData_1(wireIn[181]), .outData_0(wireOut[180]), .outData_1(wireOut[181]), .ctrl(ctrl[90]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_91(.inData_0(wireIn[182]), .inData_1(wireIn[183]), .outData_0(wireOut[182]), .outData_1(wireOut[183]), .ctrl(ctrl[91]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_92(.inData_0(wireIn[184]), .inData_1(wireIn[185]), .outData_0(wireOut[184]), .outData_1(wireOut[185]), .ctrl(ctrl[92]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_93(.inData_0(wireIn[186]), .inData_1(wireIn[187]), .outData_0(wireOut[186]), .outData_1(wireOut[187]), .ctrl(ctrl[93]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_94(.inData_0(wireIn[188]), .inData_1(wireIn[189]), .outData_0(wireOut[188]), .outData_1(wireOut[189]), .ctrl(ctrl[94]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_95(.inData_0(wireIn[190]), .inData_1(wireIn[191]), .outData_0(wireOut[190]), .outData_1(wireOut[191]), .ctrl(ctrl[95]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_96(.inData_0(wireIn[192]), .inData_1(wireIn[193]), .outData_0(wireOut[192]), .outData_1(wireOut[193]), .ctrl(ctrl[96]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_97(.inData_0(wireIn[194]), .inData_1(wireIn[195]), .outData_0(wireOut[194]), .outData_1(wireOut[195]), .ctrl(ctrl[97]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_98(.inData_0(wireIn[196]), .inData_1(wireIn[197]), .outData_0(wireOut[196]), .outData_1(wireOut[197]), .ctrl(ctrl[98]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_99(.inData_0(wireIn[198]), .inData_1(wireIn[199]), .outData_0(wireOut[198]), .outData_1(wireOut[199]), .ctrl(ctrl[99]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_100(.inData_0(wireIn[200]), .inData_1(wireIn[201]), .outData_0(wireOut[200]), .outData_1(wireOut[201]), .ctrl(ctrl[100]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_101(.inData_0(wireIn[202]), .inData_1(wireIn[203]), .outData_0(wireOut[202]), .outData_1(wireOut[203]), .ctrl(ctrl[101]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_102(.inData_0(wireIn[204]), .inData_1(wireIn[205]), .outData_0(wireOut[204]), .outData_1(wireOut[205]), .ctrl(ctrl[102]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_103(.inData_0(wireIn[206]), .inData_1(wireIn[207]), .outData_0(wireOut[206]), .outData_1(wireOut[207]), .ctrl(ctrl[103]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_104(.inData_0(wireIn[208]), .inData_1(wireIn[209]), .outData_0(wireOut[208]), .outData_1(wireOut[209]), .ctrl(ctrl[104]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_105(.inData_0(wireIn[210]), .inData_1(wireIn[211]), .outData_0(wireOut[210]), .outData_1(wireOut[211]), .ctrl(ctrl[105]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_106(.inData_0(wireIn[212]), .inData_1(wireIn[213]), .outData_0(wireOut[212]), .outData_1(wireOut[213]), .ctrl(ctrl[106]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_107(.inData_0(wireIn[214]), .inData_1(wireIn[215]), .outData_0(wireOut[214]), .outData_1(wireOut[215]), .ctrl(ctrl[107]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_108(.inData_0(wireIn[216]), .inData_1(wireIn[217]), .outData_0(wireOut[216]), .outData_1(wireOut[217]), .ctrl(ctrl[108]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_109(.inData_0(wireIn[218]), .inData_1(wireIn[219]), .outData_0(wireOut[218]), .outData_1(wireOut[219]), .ctrl(ctrl[109]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_110(.inData_0(wireIn[220]), .inData_1(wireIn[221]), .outData_0(wireOut[220]), .outData_1(wireOut[221]), .ctrl(ctrl[110]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_111(.inData_0(wireIn[222]), .inData_1(wireIn[223]), .outData_0(wireOut[222]), .outData_1(wireOut[223]), .ctrl(ctrl[111]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_112(.inData_0(wireIn[224]), .inData_1(wireIn[225]), .outData_0(wireOut[224]), .outData_1(wireOut[225]), .ctrl(ctrl[112]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_113(.inData_0(wireIn[226]), .inData_1(wireIn[227]), .outData_0(wireOut[226]), .outData_1(wireOut[227]), .ctrl(ctrl[113]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_114(.inData_0(wireIn[228]), .inData_1(wireIn[229]), .outData_0(wireOut[228]), .outData_1(wireOut[229]), .ctrl(ctrl[114]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_115(.inData_0(wireIn[230]), .inData_1(wireIn[231]), .outData_0(wireOut[230]), .outData_1(wireOut[231]), .ctrl(ctrl[115]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_116(.inData_0(wireIn[232]), .inData_1(wireIn[233]), .outData_0(wireOut[232]), .outData_1(wireOut[233]), .ctrl(ctrl[116]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_117(.inData_0(wireIn[234]), .inData_1(wireIn[235]), .outData_0(wireOut[234]), .outData_1(wireOut[235]), .ctrl(ctrl[117]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_118(.inData_0(wireIn[236]), .inData_1(wireIn[237]), .outData_0(wireOut[236]), .outData_1(wireOut[237]), .ctrl(ctrl[118]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_119(.inData_0(wireIn[238]), .inData_1(wireIn[239]), .outData_0(wireOut[238]), .outData_1(wireOut[239]), .ctrl(ctrl[119]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_120(.inData_0(wireIn[240]), .inData_1(wireIn[241]), .outData_0(wireOut[240]), .outData_1(wireOut[241]), .ctrl(ctrl[120]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_121(.inData_0(wireIn[242]), .inData_1(wireIn[243]), .outData_0(wireOut[242]), .outData_1(wireOut[243]), .ctrl(ctrl[121]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_122(.inData_0(wireIn[244]), .inData_1(wireIn[245]), .outData_0(wireOut[244]), .outData_1(wireOut[245]), .ctrl(ctrl[122]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_123(.inData_0(wireIn[246]), .inData_1(wireIn[247]), .outData_0(wireOut[246]), .outData_1(wireOut[247]), .ctrl(ctrl[123]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_124(.inData_0(wireIn[248]), .inData_1(wireIn[249]), .outData_0(wireOut[248]), .outData_1(wireOut[249]), .ctrl(ctrl[124]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_125(.inData_0(wireIn[250]), .inData_1(wireIn[251]), .outData_0(wireOut[250]), .outData_1(wireOut[251]), .ctrl(ctrl[125]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_126(.inData_0(wireIn[252]), .inData_1(wireIn[253]), .outData_0(wireOut[252]), .outData_1(wireOut[253]), .ctrl(ctrl[126]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_127(.inData_0(wireIn[254]), .inData_1(wireIn[255]), .outData_0(wireOut[254]), .outData_1(wireOut[255]), .ctrl(ctrl[127]), .clk(clk), .rst(rst));
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module wireCon_dp256_st1_L(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  assign wireOut[0] = wireIn[0];    
  assign wireOut[1] = wireIn[2];    
  assign wireOut[2] = wireIn[4];    
  assign wireOut[3] = wireIn[6];    
  assign wireOut[4] = wireIn[8];    
  assign wireOut[5] = wireIn[10];    
  assign wireOut[6] = wireIn[12];    
  assign wireOut[7] = wireIn[14];    
  assign wireOut[8] = wireIn[16];    
  assign wireOut[9] = wireIn[18];    
  assign wireOut[10] = wireIn[20];    
  assign wireOut[11] = wireIn[22];    
  assign wireOut[12] = wireIn[24];    
  assign wireOut[13] = wireIn[26];    
  assign wireOut[14] = wireIn[28];    
  assign wireOut[15] = wireIn[30];    
  assign wireOut[16] = wireIn[32];    
  assign wireOut[17] = wireIn[34];    
  assign wireOut[18] = wireIn[36];    
  assign wireOut[19] = wireIn[38];    
  assign wireOut[20] = wireIn[40];    
  assign wireOut[21] = wireIn[42];    
  assign wireOut[22] = wireIn[44];    
  assign wireOut[23] = wireIn[46];    
  assign wireOut[24] = wireIn[48];    
  assign wireOut[25] = wireIn[50];    
  assign wireOut[26] = wireIn[52];    
  assign wireOut[27] = wireIn[54];    
  assign wireOut[28] = wireIn[56];    
  assign wireOut[29] = wireIn[58];    
  assign wireOut[30] = wireIn[60];    
  assign wireOut[31] = wireIn[62];    
  assign wireOut[32] = wireIn[64];    
  assign wireOut[33] = wireIn[66];    
  assign wireOut[34] = wireIn[68];    
  assign wireOut[35] = wireIn[70];    
  assign wireOut[36] = wireIn[72];    
  assign wireOut[37] = wireIn[74];    
  assign wireOut[38] = wireIn[76];    
  assign wireOut[39] = wireIn[78];    
  assign wireOut[40] = wireIn[80];    
  assign wireOut[41] = wireIn[82];    
  assign wireOut[42] = wireIn[84];    
  assign wireOut[43] = wireIn[86];    
  assign wireOut[44] = wireIn[88];    
  assign wireOut[45] = wireIn[90];    
  assign wireOut[46] = wireIn[92];    
  assign wireOut[47] = wireIn[94];    
  assign wireOut[48] = wireIn[96];    
  assign wireOut[49] = wireIn[98];    
  assign wireOut[50] = wireIn[100];    
  assign wireOut[51] = wireIn[102];    
  assign wireOut[52] = wireIn[104];    
  assign wireOut[53] = wireIn[106];    
  assign wireOut[54] = wireIn[108];    
  assign wireOut[55] = wireIn[110];    
  assign wireOut[56] = wireIn[112];    
  assign wireOut[57] = wireIn[114];    
  assign wireOut[58] = wireIn[116];    
  assign wireOut[59] = wireIn[118];    
  assign wireOut[60] = wireIn[120];    
  assign wireOut[61] = wireIn[122];    
  assign wireOut[62] = wireIn[124];    
  assign wireOut[63] = wireIn[126];    
  assign wireOut[64] = wireIn[1];    
  assign wireOut[65] = wireIn[3];    
  assign wireOut[66] = wireIn[5];    
  assign wireOut[67] = wireIn[7];    
  assign wireOut[68] = wireIn[9];    
  assign wireOut[69] = wireIn[11];    
  assign wireOut[70] = wireIn[13];    
  assign wireOut[71] = wireIn[15];    
  assign wireOut[72] = wireIn[17];    
  assign wireOut[73] = wireIn[19];    
  assign wireOut[74] = wireIn[21];    
  assign wireOut[75] = wireIn[23];    
  assign wireOut[76] = wireIn[25];    
  assign wireOut[77] = wireIn[27];    
  assign wireOut[78] = wireIn[29];    
  assign wireOut[79] = wireIn[31];    
  assign wireOut[80] = wireIn[33];    
  assign wireOut[81] = wireIn[35];    
  assign wireOut[82] = wireIn[37];    
  assign wireOut[83] = wireIn[39];    
  assign wireOut[84] = wireIn[41];    
  assign wireOut[85] = wireIn[43];    
  assign wireOut[86] = wireIn[45];    
  assign wireOut[87] = wireIn[47];    
  assign wireOut[88] = wireIn[49];    
  assign wireOut[89] = wireIn[51];    
  assign wireOut[90] = wireIn[53];    
  assign wireOut[91] = wireIn[55];    
  assign wireOut[92] = wireIn[57];    
  assign wireOut[93] = wireIn[59];    
  assign wireOut[94] = wireIn[61];    
  assign wireOut[95] = wireIn[63];    
  assign wireOut[96] = wireIn[65];    
  assign wireOut[97] = wireIn[67];    
  assign wireOut[98] = wireIn[69];    
  assign wireOut[99] = wireIn[71];    
  assign wireOut[100] = wireIn[73];    
  assign wireOut[101] = wireIn[75];    
  assign wireOut[102] = wireIn[77];    
  assign wireOut[103] = wireIn[79];    
  assign wireOut[104] = wireIn[81];    
  assign wireOut[105] = wireIn[83];    
  assign wireOut[106] = wireIn[85];    
  assign wireOut[107] = wireIn[87];    
  assign wireOut[108] = wireIn[89];    
  assign wireOut[109] = wireIn[91];    
  assign wireOut[110] = wireIn[93];    
  assign wireOut[111] = wireIn[95];    
  assign wireOut[112] = wireIn[97];    
  assign wireOut[113] = wireIn[99];    
  assign wireOut[114] = wireIn[101];    
  assign wireOut[115] = wireIn[103];    
  assign wireOut[116] = wireIn[105];    
  assign wireOut[117] = wireIn[107];    
  assign wireOut[118] = wireIn[109];    
  assign wireOut[119] = wireIn[111];    
  assign wireOut[120] = wireIn[113];    
  assign wireOut[121] = wireIn[115];    
  assign wireOut[122] = wireIn[117];    
  assign wireOut[123] = wireIn[119];    
  assign wireOut[124] = wireIn[121];    
  assign wireOut[125] = wireIn[123];    
  assign wireOut[126] = wireIn[125];    
  assign wireOut[127] = wireIn[127];    
  assign wireOut[128] = wireIn[128];    
  assign wireOut[129] = wireIn[130];    
  assign wireOut[130] = wireIn[132];    
  assign wireOut[131] = wireIn[134];    
  assign wireOut[132] = wireIn[136];    
  assign wireOut[133] = wireIn[138];    
  assign wireOut[134] = wireIn[140];    
  assign wireOut[135] = wireIn[142];    
  assign wireOut[136] = wireIn[144];    
  assign wireOut[137] = wireIn[146];    
  assign wireOut[138] = wireIn[148];    
  assign wireOut[139] = wireIn[150];    
  assign wireOut[140] = wireIn[152];    
  assign wireOut[141] = wireIn[154];    
  assign wireOut[142] = wireIn[156];    
  assign wireOut[143] = wireIn[158];    
  assign wireOut[144] = wireIn[160];    
  assign wireOut[145] = wireIn[162];    
  assign wireOut[146] = wireIn[164];    
  assign wireOut[147] = wireIn[166];    
  assign wireOut[148] = wireIn[168];    
  assign wireOut[149] = wireIn[170];    
  assign wireOut[150] = wireIn[172];    
  assign wireOut[151] = wireIn[174];    
  assign wireOut[152] = wireIn[176];    
  assign wireOut[153] = wireIn[178];    
  assign wireOut[154] = wireIn[180];    
  assign wireOut[155] = wireIn[182];    
  assign wireOut[156] = wireIn[184];    
  assign wireOut[157] = wireIn[186];    
  assign wireOut[158] = wireIn[188];    
  assign wireOut[159] = wireIn[190];    
  assign wireOut[160] = wireIn[192];    
  assign wireOut[161] = wireIn[194];    
  assign wireOut[162] = wireIn[196];    
  assign wireOut[163] = wireIn[198];    
  assign wireOut[164] = wireIn[200];    
  assign wireOut[165] = wireIn[202];    
  assign wireOut[166] = wireIn[204];    
  assign wireOut[167] = wireIn[206];    
  assign wireOut[168] = wireIn[208];    
  assign wireOut[169] = wireIn[210];    
  assign wireOut[170] = wireIn[212];    
  assign wireOut[171] = wireIn[214];    
  assign wireOut[172] = wireIn[216];    
  assign wireOut[173] = wireIn[218];    
  assign wireOut[174] = wireIn[220];    
  assign wireOut[175] = wireIn[222];    
  assign wireOut[176] = wireIn[224];    
  assign wireOut[177] = wireIn[226];    
  assign wireOut[178] = wireIn[228];    
  assign wireOut[179] = wireIn[230];    
  assign wireOut[180] = wireIn[232];    
  assign wireOut[181] = wireIn[234];    
  assign wireOut[182] = wireIn[236];    
  assign wireOut[183] = wireIn[238];    
  assign wireOut[184] = wireIn[240];    
  assign wireOut[185] = wireIn[242];    
  assign wireOut[186] = wireIn[244];    
  assign wireOut[187] = wireIn[246];    
  assign wireOut[188] = wireIn[248];    
  assign wireOut[189] = wireIn[250];    
  assign wireOut[190] = wireIn[252];    
  assign wireOut[191] = wireIn[254];    
  assign wireOut[192] = wireIn[129];    
  assign wireOut[193] = wireIn[131];    
  assign wireOut[194] = wireIn[133];    
  assign wireOut[195] = wireIn[135];    
  assign wireOut[196] = wireIn[137];    
  assign wireOut[197] = wireIn[139];    
  assign wireOut[198] = wireIn[141];    
  assign wireOut[199] = wireIn[143];    
  assign wireOut[200] = wireIn[145];    
  assign wireOut[201] = wireIn[147];    
  assign wireOut[202] = wireIn[149];    
  assign wireOut[203] = wireIn[151];    
  assign wireOut[204] = wireIn[153];    
  assign wireOut[205] = wireIn[155];    
  assign wireOut[206] = wireIn[157];    
  assign wireOut[207] = wireIn[159];    
  assign wireOut[208] = wireIn[161];    
  assign wireOut[209] = wireIn[163];    
  assign wireOut[210] = wireIn[165];    
  assign wireOut[211] = wireIn[167];    
  assign wireOut[212] = wireIn[169];    
  assign wireOut[213] = wireIn[171];    
  assign wireOut[214] = wireIn[173];    
  assign wireOut[215] = wireIn[175];    
  assign wireOut[216] = wireIn[177];    
  assign wireOut[217] = wireIn[179];    
  assign wireOut[218] = wireIn[181];    
  assign wireOut[219] = wireIn[183];    
  assign wireOut[220] = wireIn[185];    
  assign wireOut[221] = wireIn[187];    
  assign wireOut[222] = wireIn[189];    
  assign wireOut[223] = wireIn[191];    
  assign wireOut[224] = wireIn[193];    
  assign wireOut[225] = wireIn[195];    
  assign wireOut[226] = wireIn[197];    
  assign wireOut[227] = wireIn[199];    
  assign wireOut[228] = wireIn[201];    
  assign wireOut[229] = wireIn[203];    
  assign wireOut[230] = wireIn[205];    
  assign wireOut[231] = wireIn[207];    
  assign wireOut[232] = wireIn[209];    
  assign wireOut[233] = wireIn[211];    
  assign wireOut[234] = wireIn[213];    
  assign wireOut[235] = wireIn[215];    
  assign wireOut[236] = wireIn[217];    
  assign wireOut[237] = wireIn[219];    
  assign wireOut[238] = wireIn[221];    
  assign wireOut[239] = wireIn[223];    
  assign wireOut[240] = wireIn[225];    
  assign wireOut[241] = wireIn[227];    
  assign wireOut[242] = wireIn[229];    
  assign wireOut[243] = wireIn[231];    
  assign wireOut[244] = wireIn[233];    
  assign wireOut[245] = wireIn[235];    
  assign wireOut[246] = wireIn[237];    
  assign wireOut[247] = wireIn[239];    
  assign wireOut[248] = wireIn[241];    
  assign wireOut[249] = wireIn[243];    
  assign wireOut[250] = wireIn[245];    
  assign wireOut[251] = wireIn[247];    
  assign wireOut[252] = wireIn[249];    
  assign wireOut[253] = wireIn[251];    
  assign wireOut[254] = wireIn[253];    
  assign wireOut[255] = wireIn[255];    
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module switches_stage_st2_0_L(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
ctrl,                            
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;                   
  input [128-1:0] ctrl;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  switch_2_2 switch_inst_0(.inData_0(wireIn[0]), .inData_1(wireIn[1]), .outData_0(wireOut[0]), .outData_1(wireOut[1]), .ctrl(ctrl[0]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_1(.inData_0(wireIn[2]), .inData_1(wireIn[3]), .outData_0(wireOut[2]), .outData_1(wireOut[3]), .ctrl(ctrl[1]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_2(.inData_0(wireIn[4]), .inData_1(wireIn[5]), .outData_0(wireOut[4]), .outData_1(wireOut[5]), .ctrl(ctrl[2]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_3(.inData_0(wireIn[6]), .inData_1(wireIn[7]), .outData_0(wireOut[6]), .outData_1(wireOut[7]), .ctrl(ctrl[3]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_4(.inData_0(wireIn[8]), .inData_1(wireIn[9]), .outData_0(wireOut[8]), .outData_1(wireOut[9]), .ctrl(ctrl[4]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_5(.inData_0(wireIn[10]), .inData_1(wireIn[11]), .outData_0(wireOut[10]), .outData_1(wireOut[11]), .ctrl(ctrl[5]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_6(.inData_0(wireIn[12]), .inData_1(wireIn[13]), .outData_0(wireOut[12]), .outData_1(wireOut[13]), .ctrl(ctrl[6]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_7(.inData_0(wireIn[14]), .inData_1(wireIn[15]), .outData_0(wireOut[14]), .outData_1(wireOut[15]), .ctrl(ctrl[7]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_8(.inData_0(wireIn[16]), .inData_1(wireIn[17]), .outData_0(wireOut[16]), .outData_1(wireOut[17]), .ctrl(ctrl[8]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_9(.inData_0(wireIn[18]), .inData_1(wireIn[19]), .outData_0(wireOut[18]), .outData_1(wireOut[19]), .ctrl(ctrl[9]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_10(.inData_0(wireIn[20]), .inData_1(wireIn[21]), .outData_0(wireOut[20]), .outData_1(wireOut[21]), .ctrl(ctrl[10]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_11(.inData_0(wireIn[22]), .inData_1(wireIn[23]), .outData_0(wireOut[22]), .outData_1(wireOut[23]), .ctrl(ctrl[11]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_12(.inData_0(wireIn[24]), .inData_1(wireIn[25]), .outData_0(wireOut[24]), .outData_1(wireOut[25]), .ctrl(ctrl[12]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_13(.inData_0(wireIn[26]), .inData_1(wireIn[27]), .outData_0(wireOut[26]), .outData_1(wireOut[27]), .ctrl(ctrl[13]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_14(.inData_0(wireIn[28]), .inData_1(wireIn[29]), .outData_0(wireOut[28]), .outData_1(wireOut[29]), .ctrl(ctrl[14]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_15(.inData_0(wireIn[30]), .inData_1(wireIn[31]), .outData_0(wireOut[30]), .outData_1(wireOut[31]), .ctrl(ctrl[15]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_16(.inData_0(wireIn[32]), .inData_1(wireIn[33]), .outData_0(wireOut[32]), .outData_1(wireOut[33]), .ctrl(ctrl[16]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_17(.inData_0(wireIn[34]), .inData_1(wireIn[35]), .outData_0(wireOut[34]), .outData_1(wireOut[35]), .ctrl(ctrl[17]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_18(.inData_0(wireIn[36]), .inData_1(wireIn[37]), .outData_0(wireOut[36]), .outData_1(wireOut[37]), .ctrl(ctrl[18]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_19(.inData_0(wireIn[38]), .inData_1(wireIn[39]), .outData_0(wireOut[38]), .outData_1(wireOut[39]), .ctrl(ctrl[19]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_20(.inData_0(wireIn[40]), .inData_1(wireIn[41]), .outData_0(wireOut[40]), .outData_1(wireOut[41]), .ctrl(ctrl[20]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_21(.inData_0(wireIn[42]), .inData_1(wireIn[43]), .outData_0(wireOut[42]), .outData_1(wireOut[43]), .ctrl(ctrl[21]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_22(.inData_0(wireIn[44]), .inData_1(wireIn[45]), .outData_0(wireOut[44]), .outData_1(wireOut[45]), .ctrl(ctrl[22]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_23(.inData_0(wireIn[46]), .inData_1(wireIn[47]), .outData_0(wireOut[46]), .outData_1(wireOut[47]), .ctrl(ctrl[23]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_24(.inData_0(wireIn[48]), .inData_1(wireIn[49]), .outData_0(wireOut[48]), .outData_1(wireOut[49]), .ctrl(ctrl[24]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_25(.inData_0(wireIn[50]), .inData_1(wireIn[51]), .outData_0(wireOut[50]), .outData_1(wireOut[51]), .ctrl(ctrl[25]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_26(.inData_0(wireIn[52]), .inData_1(wireIn[53]), .outData_0(wireOut[52]), .outData_1(wireOut[53]), .ctrl(ctrl[26]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_27(.inData_0(wireIn[54]), .inData_1(wireIn[55]), .outData_0(wireOut[54]), .outData_1(wireOut[55]), .ctrl(ctrl[27]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_28(.inData_0(wireIn[56]), .inData_1(wireIn[57]), .outData_0(wireOut[56]), .outData_1(wireOut[57]), .ctrl(ctrl[28]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_29(.inData_0(wireIn[58]), .inData_1(wireIn[59]), .outData_0(wireOut[58]), .outData_1(wireOut[59]), .ctrl(ctrl[29]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_30(.inData_0(wireIn[60]), .inData_1(wireIn[61]), .outData_0(wireOut[60]), .outData_1(wireOut[61]), .ctrl(ctrl[30]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_31(.inData_0(wireIn[62]), .inData_1(wireIn[63]), .outData_0(wireOut[62]), .outData_1(wireOut[63]), .ctrl(ctrl[31]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_32(.inData_0(wireIn[64]), .inData_1(wireIn[65]), .outData_0(wireOut[64]), .outData_1(wireOut[65]), .ctrl(ctrl[32]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_33(.inData_0(wireIn[66]), .inData_1(wireIn[67]), .outData_0(wireOut[66]), .outData_1(wireOut[67]), .ctrl(ctrl[33]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_34(.inData_0(wireIn[68]), .inData_1(wireIn[69]), .outData_0(wireOut[68]), .outData_1(wireOut[69]), .ctrl(ctrl[34]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_35(.inData_0(wireIn[70]), .inData_1(wireIn[71]), .outData_0(wireOut[70]), .outData_1(wireOut[71]), .ctrl(ctrl[35]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_36(.inData_0(wireIn[72]), .inData_1(wireIn[73]), .outData_0(wireOut[72]), .outData_1(wireOut[73]), .ctrl(ctrl[36]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_37(.inData_0(wireIn[74]), .inData_1(wireIn[75]), .outData_0(wireOut[74]), .outData_1(wireOut[75]), .ctrl(ctrl[37]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_38(.inData_0(wireIn[76]), .inData_1(wireIn[77]), .outData_0(wireOut[76]), .outData_1(wireOut[77]), .ctrl(ctrl[38]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_39(.inData_0(wireIn[78]), .inData_1(wireIn[79]), .outData_0(wireOut[78]), .outData_1(wireOut[79]), .ctrl(ctrl[39]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_40(.inData_0(wireIn[80]), .inData_1(wireIn[81]), .outData_0(wireOut[80]), .outData_1(wireOut[81]), .ctrl(ctrl[40]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_41(.inData_0(wireIn[82]), .inData_1(wireIn[83]), .outData_0(wireOut[82]), .outData_1(wireOut[83]), .ctrl(ctrl[41]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_42(.inData_0(wireIn[84]), .inData_1(wireIn[85]), .outData_0(wireOut[84]), .outData_1(wireOut[85]), .ctrl(ctrl[42]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_43(.inData_0(wireIn[86]), .inData_1(wireIn[87]), .outData_0(wireOut[86]), .outData_1(wireOut[87]), .ctrl(ctrl[43]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_44(.inData_0(wireIn[88]), .inData_1(wireIn[89]), .outData_0(wireOut[88]), .outData_1(wireOut[89]), .ctrl(ctrl[44]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_45(.inData_0(wireIn[90]), .inData_1(wireIn[91]), .outData_0(wireOut[90]), .outData_1(wireOut[91]), .ctrl(ctrl[45]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_46(.inData_0(wireIn[92]), .inData_1(wireIn[93]), .outData_0(wireOut[92]), .outData_1(wireOut[93]), .ctrl(ctrl[46]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_47(.inData_0(wireIn[94]), .inData_1(wireIn[95]), .outData_0(wireOut[94]), .outData_1(wireOut[95]), .ctrl(ctrl[47]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_48(.inData_0(wireIn[96]), .inData_1(wireIn[97]), .outData_0(wireOut[96]), .outData_1(wireOut[97]), .ctrl(ctrl[48]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_49(.inData_0(wireIn[98]), .inData_1(wireIn[99]), .outData_0(wireOut[98]), .outData_1(wireOut[99]), .ctrl(ctrl[49]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_50(.inData_0(wireIn[100]), .inData_1(wireIn[101]), .outData_0(wireOut[100]), .outData_1(wireOut[101]), .ctrl(ctrl[50]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_51(.inData_0(wireIn[102]), .inData_1(wireIn[103]), .outData_0(wireOut[102]), .outData_1(wireOut[103]), .ctrl(ctrl[51]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_52(.inData_0(wireIn[104]), .inData_1(wireIn[105]), .outData_0(wireOut[104]), .outData_1(wireOut[105]), .ctrl(ctrl[52]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_53(.inData_0(wireIn[106]), .inData_1(wireIn[107]), .outData_0(wireOut[106]), .outData_1(wireOut[107]), .ctrl(ctrl[53]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_54(.inData_0(wireIn[108]), .inData_1(wireIn[109]), .outData_0(wireOut[108]), .outData_1(wireOut[109]), .ctrl(ctrl[54]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_55(.inData_0(wireIn[110]), .inData_1(wireIn[111]), .outData_0(wireOut[110]), .outData_1(wireOut[111]), .ctrl(ctrl[55]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_56(.inData_0(wireIn[112]), .inData_1(wireIn[113]), .outData_0(wireOut[112]), .outData_1(wireOut[113]), .ctrl(ctrl[56]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_57(.inData_0(wireIn[114]), .inData_1(wireIn[115]), .outData_0(wireOut[114]), .outData_1(wireOut[115]), .ctrl(ctrl[57]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_58(.inData_0(wireIn[116]), .inData_1(wireIn[117]), .outData_0(wireOut[116]), .outData_1(wireOut[117]), .ctrl(ctrl[58]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_59(.inData_0(wireIn[118]), .inData_1(wireIn[119]), .outData_0(wireOut[118]), .outData_1(wireOut[119]), .ctrl(ctrl[59]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_60(.inData_0(wireIn[120]), .inData_1(wireIn[121]), .outData_0(wireOut[120]), .outData_1(wireOut[121]), .ctrl(ctrl[60]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_61(.inData_0(wireIn[122]), .inData_1(wireIn[123]), .outData_0(wireOut[122]), .outData_1(wireOut[123]), .ctrl(ctrl[61]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_62(.inData_0(wireIn[124]), .inData_1(wireIn[125]), .outData_0(wireOut[124]), .outData_1(wireOut[125]), .ctrl(ctrl[62]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_63(.inData_0(wireIn[126]), .inData_1(wireIn[127]), .outData_0(wireOut[126]), .outData_1(wireOut[127]), .ctrl(ctrl[63]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_64(.inData_0(wireIn[128]), .inData_1(wireIn[129]), .outData_0(wireOut[128]), .outData_1(wireOut[129]), .ctrl(ctrl[64]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_65(.inData_0(wireIn[130]), .inData_1(wireIn[131]), .outData_0(wireOut[130]), .outData_1(wireOut[131]), .ctrl(ctrl[65]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_66(.inData_0(wireIn[132]), .inData_1(wireIn[133]), .outData_0(wireOut[132]), .outData_1(wireOut[133]), .ctrl(ctrl[66]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_67(.inData_0(wireIn[134]), .inData_1(wireIn[135]), .outData_0(wireOut[134]), .outData_1(wireOut[135]), .ctrl(ctrl[67]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_68(.inData_0(wireIn[136]), .inData_1(wireIn[137]), .outData_0(wireOut[136]), .outData_1(wireOut[137]), .ctrl(ctrl[68]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_69(.inData_0(wireIn[138]), .inData_1(wireIn[139]), .outData_0(wireOut[138]), .outData_1(wireOut[139]), .ctrl(ctrl[69]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_70(.inData_0(wireIn[140]), .inData_1(wireIn[141]), .outData_0(wireOut[140]), .outData_1(wireOut[141]), .ctrl(ctrl[70]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_71(.inData_0(wireIn[142]), .inData_1(wireIn[143]), .outData_0(wireOut[142]), .outData_1(wireOut[143]), .ctrl(ctrl[71]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_72(.inData_0(wireIn[144]), .inData_1(wireIn[145]), .outData_0(wireOut[144]), .outData_1(wireOut[145]), .ctrl(ctrl[72]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_73(.inData_0(wireIn[146]), .inData_1(wireIn[147]), .outData_0(wireOut[146]), .outData_1(wireOut[147]), .ctrl(ctrl[73]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_74(.inData_0(wireIn[148]), .inData_1(wireIn[149]), .outData_0(wireOut[148]), .outData_1(wireOut[149]), .ctrl(ctrl[74]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_75(.inData_0(wireIn[150]), .inData_1(wireIn[151]), .outData_0(wireOut[150]), .outData_1(wireOut[151]), .ctrl(ctrl[75]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_76(.inData_0(wireIn[152]), .inData_1(wireIn[153]), .outData_0(wireOut[152]), .outData_1(wireOut[153]), .ctrl(ctrl[76]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_77(.inData_0(wireIn[154]), .inData_1(wireIn[155]), .outData_0(wireOut[154]), .outData_1(wireOut[155]), .ctrl(ctrl[77]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_78(.inData_0(wireIn[156]), .inData_1(wireIn[157]), .outData_0(wireOut[156]), .outData_1(wireOut[157]), .ctrl(ctrl[78]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_79(.inData_0(wireIn[158]), .inData_1(wireIn[159]), .outData_0(wireOut[158]), .outData_1(wireOut[159]), .ctrl(ctrl[79]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_80(.inData_0(wireIn[160]), .inData_1(wireIn[161]), .outData_0(wireOut[160]), .outData_1(wireOut[161]), .ctrl(ctrl[80]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_81(.inData_0(wireIn[162]), .inData_1(wireIn[163]), .outData_0(wireOut[162]), .outData_1(wireOut[163]), .ctrl(ctrl[81]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_82(.inData_0(wireIn[164]), .inData_1(wireIn[165]), .outData_0(wireOut[164]), .outData_1(wireOut[165]), .ctrl(ctrl[82]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_83(.inData_0(wireIn[166]), .inData_1(wireIn[167]), .outData_0(wireOut[166]), .outData_1(wireOut[167]), .ctrl(ctrl[83]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_84(.inData_0(wireIn[168]), .inData_1(wireIn[169]), .outData_0(wireOut[168]), .outData_1(wireOut[169]), .ctrl(ctrl[84]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_85(.inData_0(wireIn[170]), .inData_1(wireIn[171]), .outData_0(wireOut[170]), .outData_1(wireOut[171]), .ctrl(ctrl[85]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_86(.inData_0(wireIn[172]), .inData_1(wireIn[173]), .outData_0(wireOut[172]), .outData_1(wireOut[173]), .ctrl(ctrl[86]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_87(.inData_0(wireIn[174]), .inData_1(wireIn[175]), .outData_0(wireOut[174]), .outData_1(wireOut[175]), .ctrl(ctrl[87]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_88(.inData_0(wireIn[176]), .inData_1(wireIn[177]), .outData_0(wireOut[176]), .outData_1(wireOut[177]), .ctrl(ctrl[88]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_89(.inData_0(wireIn[178]), .inData_1(wireIn[179]), .outData_0(wireOut[178]), .outData_1(wireOut[179]), .ctrl(ctrl[89]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_90(.inData_0(wireIn[180]), .inData_1(wireIn[181]), .outData_0(wireOut[180]), .outData_1(wireOut[181]), .ctrl(ctrl[90]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_91(.inData_0(wireIn[182]), .inData_1(wireIn[183]), .outData_0(wireOut[182]), .outData_1(wireOut[183]), .ctrl(ctrl[91]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_92(.inData_0(wireIn[184]), .inData_1(wireIn[185]), .outData_0(wireOut[184]), .outData_1(wireOut[185]), .ctrl(ctrl[92]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_93(.inData_0(wireIn[186]), .inData_1(wireIn[187]), .outData_0(wireOut[186]), .outData_1(wireOut[187]), .ctrl(ctrl[93]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_94(.inData_0(wireIn[188]), .inData_1(wireIn[189]), .outData_0(wireOut[188]), .outData_1(wireOut[189]), .ctrl(ctrl[94]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_95(.inData_0(wireIn[190]), .inData_1(wireIn[191]), .outData_0(wireOut[190]), .outData_1(wireOut[191]), .ctrl(ctrl[95]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_96(.inData_0(wireIn[192]), .inData_1(wireIn[193]), .outData_0(wireOut[192]), .outData_1(wireOut[193]), .ctrl(ctrl[96]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_97(.inData_0(wireIn[194]), .inData_1(wireIn[195]), .outData_0(wireOut[194]), .outData_1(wireOut[195]), .ctrl(ctrl[97]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_98(.inData_0(wireIn[196]), .inData_1(wireIn[197]), .outData_0(wireOut[196]), .outData_1(wireOut[197]), .ctrl(ctrl[98]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_99(.inData_0(wireIn[198]), .inData_1(wireIn[199]), .outData_0(wireOut[198]), .outData_1(wireOut[199]), .ctrl(ctrl[99]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_100(.inData_0(wireIn[200]), .inData_1(wireIn[201]), .outData_0(wireOut[200]), .outData_1(wireOut[201]), .ctrl(ctrl[100]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_101(.inData_0(wireIn[202]), .inData_1(wireIn[203]), .outData_0(wireOut[202]), .outData_1(wireOut[203]), .ctrl(ctrl[101]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_102(.inData_0(wireIn[204]), .inData_1(wireIn[205]), .outData_0(wireOut[204]), .outData_1(wireOut[205]), .ctrl(ctrl[102]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_103(.inData_0(wireIn[206]), .inData_1(wireIn[207]), .outData_0(wireOut[206]), .outData_1(wireOut[207]), .ctrl(ctrl[103]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_104(.inData_0(wireIn[208]), .inData_1(wireIn[209]), .outData_0(wireOut[208]), .outData_1(wireOut[209]), .ctrl(ctrl[104]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_105(.inData_0(wireIn[210]), .inData_1(wireIn[211]), .outData_0(wireOut[210]), .outData_1(wireOut[211]), .ctrl(ctrl[105]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_106(.inData_0(wireIn[212]), .inData_1(wireIn[213]), .outData_0(wireOut[212]), .outData_1(wireOut[213]), .ctrl(ctrl[106]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_107(.inData_0(wireIn[214]), .inData_1(wireIn[215]), .outData_0(wireOut[214]), .outData_1(wireOut[215]), .ctrl(ctrl[107]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_108(.inData_0(wireIn[216]), .inData_1(wireIn[217]), .outData_0(wireOut[216]), .outData_1(wireOut[217]), .ctrl(ctrl[108]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_109(.inData_0(wireIn[218]), .inData_1(wireIn[219]), .outData_0(wireOut[218]), .outData_1(wireOut[219]), .ctrl(ctrl[109]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_110(.inData_0(wireIn[220]), .inData_1(wireIn[221]), .outData_0(wireOut[220]), .outData_1(wireOut[221]), .ctrl(ctrl[110]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_111(.inData_0(wireIn[222]), .inData_1(wireIn[223]), .outData_0(wireOut[222]), .outData_1(wireOut[223]), .ctrl(ctrl[111]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_112(.inData_0(wireIn[224]), .inData_1(wireIn[225]), .outData_0(wireOut[224]), .outData_1(wireOut[225]), .ctrl(ctrl[112]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_113(.inData_0(wireIn[226]), .inData_1(wireIn[227]), .outData_0(wireOut[226]), .outData_1(wireOut[227]), .ctrl(ctrl[113]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_114(.inData_0(wireIn[228]), .inData_1(wireIn[229]), .outData_0(wireOut[228]), .outData_1(wireOut[229]), .ctrl(ctrl[114]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_115(.inData_0(wireIn[230]), .inData_1(wireIn[231]), .outData_0(wireOut[230]), .outData_1(wireOut[231]), .ctrl(ctrl[115]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_116(.inData_0(wireIn[232]), .inData_1(wireIn[233]), .outData_0(wireOut[232]), .outData_1(wireOut[233]), .ctrl(ctrl[116]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_117(.inData_0(wireIn[234]), .inData_1(wireIn[235]), .outData_0(wireOut[234]), .outData_1(wireOut[235]), .ctrl(ctrl[117]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_118(.inData_0(wireIn[236]), .inData_1(wireIn[237]), .outData_0(wireOut[236]), .outData_1(wireOut[237]), .ctrl(ctrl[118]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_119(.inData_0(wireIn[238]), .inData_1(wireIn[239]), .outData_0(wireOut[238]), .outData_1(wireOut[239]), .ctrl(ctrl[119]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_120(.inData_0(wireIn[240]), .inData_1(wireIn[241]), .outData_0(wireOut[240]), .outData_1(wireOut[241]), .ctrl(ctrl[120]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_121(.inData_0(wireIn[242]), .inData_1(wireIn[243]), .outData_0(wireOut[242]), .outData_1(wireOut[243]), .ctrl(ctrl[121]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_122(.inData_0(wireIn[244]), .inData_1(wireIn[245]), .outData_0(wireOut[244]), .outData_1(wireOut[245]), .ctrl(ctrl[122]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_123(.inData_0(wireIn[246]), .inData_1(wireIn[247]), .outData_0(wireOut[246]), .outData_1(wireOut[247]), .ctrl(ctrl[123]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_124(.inData_0(wireIn[248]), .inData_1(wireIn[249]), .outData_0(wireOut[248]), .outData_1(wireOut[249]), .ctrl(ctrl[124]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_125(.inData_0(wireIn[250]), .inData_1(wireIn[251]), .outData_0(wireOut[250]), .outData_1(wireOut[251]), .ctrl(ctrl[125]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_126(.inData_0(wireIn[252]), .inData_1(wireIn[253]), .outData_0(wireOut[252]), .outData_1(wireOut[253]), .ctrl(ctrl[126]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_127(.inData_0(wireIn[254]), .inData_1(wireIn[255]), .outData_0(wireOut[254]), .outData_1(wireOut[255]), .ctrl(ctrl[127]), .clk(clk), .rst(rst));
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module wireCon_dp256_st2_L(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  assign wireOut[0] = wireIn[0];    
  assign wireOut[1] = wireIn[2];    
  assign wireOut[2] = wireIn[4];    
  assign wireOut[3] = wireIn[6];    
  assign wireOut[4] = wireIn[8];    
  assign wireOut[5] = wireIn[10];    
  assign wireOut[6] = wireIn[12];    
  assign wireOut[7] = wireIn[14];    
  assign wireOut[8] = wireIn[16];    
  assign wireOut[9] = wireIn[18];    
  assign wireOut[10] = wireIn[20];    
  assign wireOut[11] = wireIn[22];    
  assign wireOut[12] = wireIn[24];    
  assign wireOut[13] = wireIn[26];    
  assign wireOut[14] = wireIn[28];    
  assign wireOut[15] = wireIn[30];    
  assign wireOut[16] = wireIn[32];    
  assign wireOut[17] = wireIn[34];    
  assign wireOut[18] = wireIn[36];    
  assign wireOut[19] = wireIn[38];    
  assign wireOut[20] = wireIn[40];    
  assign wireOut[21] = wireIn[42];    
  assign wireOut[22] = wireIn[44];    
  assign wireOut[23] = wireIn[46];    
  assign wireOut[24] = wireIn[48];    
  assign wireOut[25] = wireIn[50];    
  assign wireOut[26] = wireIn[52];    
  assign wireOut[27] = wireIn[54];    
  assign wireOut[28] = wireIn[56];    
  assign wireOut[29] = wireIn[58];    
  assign wireOut[30] = wireIn[60];    
  assign wireOut[31] = wireIn[62];    
  assign wireOut[32] = wireIn[1];    
  assign wireOut[33] = wireIn[3];    
  assign wireOut[34] = wireIn[5];    
  assign wireOut[35] = wireIn[7];    
  assign wireOut[36] = wireIn[9];    
  assign wireOut[37] = wireIn[11];    
  assign wireOut[38] = wireIn[13];    
  assign wireOut[39] = wireIn[15];    
  assign wireOut[40] = wireIn[17];    
  assign wireOut[41] = wireIn[19];    
  assign wireOut[42] = wireIn[21];    
  assign wireOut[43] = wireIn[23];    
  assign wireOut[44] = wireIn[25];    
  assign wireOut[45] = wireIn[27];    
  assign wireOut[46] = wireIn[29];    
  assign wireOut[47] = wireIn[31];    
  assign wireOut[48] = wireIn[33];    
  assign wireOut[49] = wireIn[35];    
  assign wireOut[50] = wireIn[37];    
  assign wireOut[51] = wireIn[39];    
  assign wireOut[52] = wireIn[41];    
  assign wireOut[53] = wireIn[43];    
  assign wireOut[54] = wireIn[45];    
  assign wireOut[55] = wireIn[47];    
  assign wireOut[56] = wireIn[49];    
  assign wireOut[57] = wireIn[51];    
  assign wireOut[58] = wireIn[53];    
  assign wireOut[59] = wireIn[55];    
  assign wireOut[60] = wireIn[57];    
  assign wireOut[61] = wireIn[59];    
  assign wireOut[62] = wireIn[61];    
  assign wireOut[63] = wireIn[63];    
  assign wireOut[64] = wireIn[64];    
  assign wireOut[65] = wireIn[66];    
  assign wireOut[66] = wireIn[68];    
  assign wireOut[67] = wireIn[70];    
  assign wireOut[68] = wireIn[72];    
  assign wireOut[69] = wireIn[74];    
  assign wireOut[70] = wireIn[76];    
  assign wireOut[71] = wireIn[78];    
  assign wireOut[72] = wireIn[80];    
  assign wireOut[73] = wireIn[82];    
  assign wireOut[74] = wireIn[84];    
  assign wireOut[75] = wireIn[86];    
  assign wireOut[76] = wireIn[88];    
  assign wireOut[77] = wireIn[90];    
  assign wireOut[78] = wireIn[92];    
  assign wireOut[79] = wireIn[94];    
  assign wireOut[80] = wireIn[96];    
  assign wireOut[81] = wireIn[98];    
  assign wireOut[82] = wireIn[100];    
  assign wireOut[83] = wireIn[102];    
  assign wireOut[84] = wireIn[104];    
  assign wireOut[85] = wireIn[106];    
  assign wireOut[86] = wireIn[108];    
  assign wireOut[87] = wireIn[110];    
  assign wireOut[88] = wireIn[112];    
  assign wireOut[89] = wireIn[114];    
  assign wireOut[90] = wireIn[116];    
  assign wireOut[91] = wireIn[118];    
  assign wireOut[92] = wireIn[120];    
  assign wireOut[93] = wireIn[122];    
  assign wireOut[94] = wireIn[124];    
  assign wireOut[95] = wireIn[126];    
  assign wireOut[96] = wireIn[65];    
  assign wireOut[97] = wireIn[67];    
  assign wireOut[98] = wireIn[69];    
  assign wireOut[99] = wireIn[71];    
  assign wireOut[100] = wireIn[73];    
  assign wireOut[101] = wireIn[75];    
  assign wireOut[102] = wireIn[77];    
  assign wireOut[103] = wireIn[79];    
  assign wireOut[104] = wireIn[81];    
  assign wireOut[105] = wireIn[83];    
  assign wireOut[106] = wireIn[85];    
  assign wireOut[107] = wireIn[87];    
  assign wireOut[108] = wireIn[89];    
  assign wireOut[109] = wireIn[91];    
  assign wireOut[110] = wireIn[93];    
  assign wireOut[111] = wireIn[95];    
  assign wireOut[112] = wireIn[97];    
  assign wireOut[113] = wireIn[99];    
  assign wireOut[114] = wireIn[101];    
  assign wireOut[115] = wireIn[103];    
  assign wireOut[116] = wireIn[105];    
  assign wireOut[117] = wireIn[107];    
  assign wireOut[118] = wireIn[109];    
  assign wireOut[119] = wireIn[111];    
  assign wireOut[120] = wireIn[113];    
  assign wireOut[121] = wireIn[115];    
  assign wireOut[122] = wireIn[117];    
  assign wireOut[123] = wireIn[119];    
  assign wireOut[124] = wireIn[121];    
  assign wireOut[125] = wireIn[123];    
  assign wireOut[126] = wireIn[125];    
  assign wireOut[127] = wireIn[127];    
  assign wireOut[128] = wireIn[128];    
  assign wireOut[129] = wireIn[130];    
  assign wireOut[130] = wireIn[132];    
  assign wireOut[131] = wireIn[134];    
  assign wireOut[132] = wireIn[136];    
  assign wireOut[133] = wireIn[138];    
  assign wireOut[134] = wireIn[140];    
  assign wireOut[135] = wireIn[142];    
  assign wireOut[136] = wireIn[144];    
  assign wireOut[137] = wireIn[146];    
  assign wireOut[138] = wireIn[148];    
  assign wireOut[139] = wireIn[150];    
  assign wireOut[140] = wireIn[152];    
  assign wireOut[141] = wireIn[154];    
  assign wireOut[142] = wireIn[156];    
  assign wireOut[143] = wireIn[158];    
  assign wireOut[144] = wireIn[160];    
  assign wireOut[145] = wireIn[162];    
  assign wireOut[146] = wireIn[164];    
  assign wireOut[147] = wireIn[166];    
  assign wireOut[148] = wireIn[168];    
  assign wireOut[149] = wireIn[170];    
  assign wireOut[150] = wireIn[172];    
  assign wireOut[151] = wireIn[174];    
  assign wireOut[152] = wireIn[176];    
  assign wireOut[153] = wireIn[178];    
  assign wireOut[154] = wireIn[180];    
  assign wireOut[155] = wireIn[182];    
  assign wireOut[156] = wireIn[184];    
  assign wireOut[157] = wireIn[186];    
  assign wireOut[158] = wireIn[188];    
  assign wireOut[159] = wireIn[190];    
  assign wireOut[160] = wireIn[129];    
  assign wireOut[161] = wireIn[131];    
  assign wireOut[162] = wireIn[133];    
  assign wireOut[163] = wireIn[135];    
  assign wireOut[164] = wireIn[137];    
  assign wireOut[165] = wireIn[139];    
  assign wireOut[166] = wireIn[141];    
  assign wireOut[167] = wireIn[143];    
  assign wireOut[168] = wireIn[145];    
  assign wireOut[169] = wireIn[147];    
  assign wireOut[170] = wireIn[149];    
  assign wireOut[171] = wireIn[151];    
  assign wireOut[172] = wireIn[153];    
  assign wireOut[173] = wireIn[155];    
  assign wireOut[174] = wireIn[157];    
  assign wireOut[175] = wireIn[159];    
  assign wireOut[176] = wireIn[161];    
  assign wireOut[177] = wireIn[163];    
  assign wireOut[178] = wireIn[165];    
  assign wireOut[179] = wireIn[167];    
  assign wireOut[180] = wireIn[169];    
  assign wireOut[181] = wireIn[171];    
  assign wireOut[182] = wireIn[173];    
  assign wireOut[183] = wireIn[175];    
  assign wireOut[184] = wireIn[177];    
  assign wireOut[185] = wireIn[179];    
  assign wireOut[186] = wireIn[181];    
  assign wireOut[187] = wireIn[183];    
  assign wireOut[188] = wireIn[185];    
  assign wireOut[189] = wireIn[187];    
  assign wireOut[190] = wireIn[189];    
  assign wireOut[191] = wireIn[191];    
  assign wireOut[192] = wireIn[192];    
  assign wireOut[193] = wireIn[194];    
  assign wireOut[194] = wireIn[196];    
  assign wireOut[195] = wireIn[198];    
  assign wireOut[196] = wireIn[200];    
  assign wireOut[197] = wireIn[202];    
  assign wireOut[198] = wireIn[204];    
  assign wireOut[199] = wireIn[206];    
  assign wireOut[200] = wireIn[208];    
  assign wireOut[201] = wireIn[210];    
  assign wireOut[202] = wireIn[212];    
  assign wireOut[203] = wireIn[214];    
  assign wireOut[204] = wireIn[216];    
  assign wireOut[205] = wireIn[218];    
  assign wireOut[206] = wireIn[220];    
  assign wireOut[207] = wireIn[222];    
  assign wireOut[208] = wireIn[224];    
  assign wireOut[209] = wireIn[226];    
  assign wireOut[210] = wireIn[228];    
  assign wireOut[211] = wireIn[230];    
  assign wireOut[212] = wireIn[232];    
  assign wireOut[213] = wireIn[234];    
  assign wireOut[214] = wireIn[236];    
  assign wireOut[215] = wireIn[238];    
  assign wireOut[216] = wireIn[240];    
  assign wireOut[217] = wireIn[242];    
  assign wireOut[218] = wireIn[244];    
  assign wireOut[219] = wireIn[246];    
  assign wireOut[220] = wireIn[248];    
  assign wireOut[221] = wireIn[250];    
  assign wireOut[222] = wireIn[252];    
  assign wireOut[223] = wireIn[254];    
  assign wireOut[224] = wireIn[193];    
  assign wireOut[225] = wireIn[195];    
  assign wireOut[226] = wireIn[197];    
  assign wireOut[227] = wireIn[199];    
  assign wireOut[228] = wireIn[201];    
  assign wireOut[229] = wireIn[203];    
  assign wireOut[230] = wireIn[205];    
  assign wireOut[231] = wireIn[207];    
  assign wireOut[232] = wireIn[209];    
  assign wireOut[233] = wireIn[211];    
  assign wireOut[234] = wireIn[213];    
  assign wireOut[235] = wireIn[215];    
  assign wireOut[236] = wireIn[217];    
  assign wireOut[237] = wireIn[219];    
  assign wireOut[238] = wireIn[221];    
  assign wireOut[239] = wireIn[223];    
  assign wireOut[240] = wireIn[225];    
  assign wireOut[241] = wireIn[227];    
  assign wireOut[242] = wireIn[229];    
  assign wireOut[243] = wireIn[231];    
  assign wireOut[244] = wireIn[233];    
  assign wireOut[245] = wireIn[235];    
  assign wireOut[246] = wireIn[237];    
  assign wireOut[247] = wireIn[239];    
  assign wireOut[248] = wireIn[241];    
  assign wireOut[249] = wireIn[243];    
  assign wireOut[250] = wireIn[245];    
  assign wireOut[251] = wireIn[247];    
  assign wireOut[252] = wireIn[249];    
  assign wireOut[253] = wireIn[251];    
  assign wireOut[254] = wireIn[253];    
  assign wireOut[255] = wireIn[255];    
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module switches_stage_st3_0_L(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
ctrl,                            
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;                   
  input [128-1:0] ctrl;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  switch_2_2 switch_inst_0(.inData_0(wireIn[0]), .inData_1(wireIn[1]), .outData_0(wireOut[0]), .outData_1(wireOut[1]), .ctrl(ctrl[0]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_1(.inData_0(wireIn[2]), .inData_1(wireIn[3]), .outData_0(wireOut[2]), .outData_1(wireOut[3]), .ctrl(ctrl[1]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_2(.inData_0(wireIn[4]), .inData_1(wireIn[5]), .outData_0(wireOut[4]), .outData_1(wireOut[5]), .ctrl(ctrl[2]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_3(.inData_0(wireIn[6]), .inData_1(wireIn[7]), .outData_0(wireOut[6]), .outData_1(wireOut[7]), .ctrl(ctrl[3]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_4(.inData_0(wireIn[8]), .inData_1(wireIn[9]), .outData_0(wireOut[8]), .outData_1(wireOut[9]), .ctrl(ctrl[4]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_5(.inData_0(wireIn[10]), .inData_1(wireIn[11]), .outData_0(wireOut[10]), .outData_1(wireOut[11]), .ctrl(ctrl[5]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_6(.inData_0(wireIn[12]), .inData_1(wireIn[13]), .outData_0(wireOut[12]), .outData_1(wireOut[13]), .ctrl(ctrl[6]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_7(.inData_0(wireIn[14]), .inData_1(wireIn[15]), .outData_0(wireOut[14]), .outData_1(wireOut[15]), .ctrl(ctrl[7]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_8(.inData_0(wireIn[16]), .inData_1(wireIn[17]), .outData_0(wireOut[16]), .outData_1(wireOut[17]), .ctrl(ctrl[8]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_9(.inData_0(wireIn[18]), .inData_1(wireIn[19]), .outData_0(wireOut[18]), .outData_1(wireOut[19]), .ctrl(ctrl[9]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_10(.inData_0(wireIn[20]), .inData_1(wireIn[21]), .outData_0(wireOut[20]), .outData_1(wireOut[21]), .ctrl(ctrl[10]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_11(.inData_0(wireIn[22]), .inData_1(wireIn[23]), .outData_0(wireOut[22]), .outData_1(wireOut[23]), .ctrl(ctrl[11]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_12(.inData_0(wireIn[24]), .inData_1(wireIn[25]), .outData_0(wireOut[24]), .outData_1(wireOut[25]), .ctrl(ctrl[12]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_13(.inData_0(wireIn[26]), .inData_1(wireIn[27]), .outData_0(wireOut[26]), .outData_1(wireOut[27]), .ctrl(ctrl[13]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_14(.inData_0(wireIn[28]), .inData_1(wireIn[29]), .outData_0(wireOut[28]), .outData_1(wireOut[29]), .ctrl(ctrl[14]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_15(.inData_0(wireIn[30]), .inData_1(wireIn[31]), .outData_0(wireOut[30]), .outData_1(wireOut[31]), .ctrl(ctrl[15]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_16(.inData_0(wireIn[32]), .inData_1(wireIn[33]), .outData_0(wireOut[32]), .outData_1(wireOut[33]), .ctrl(ctrl[16]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_17(.inData_0(wireIn[34]), .inData_1(wireIn[35]), .outData_0(wireOut[34]), .outData_1(wireOut[35]), .ctrl(ctrl[17]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_18(.inData_0(wireIn[36]), .inData_1(wireIn[37]), .outData_0(wireOut[36]), .outData_1(wireOut[37]), .ctrl(ctrl[18]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_19(.inData_0(wireIn[38]), .inData_1(wireIn[39]), .outData_0(wireOut[38]), .outData_1(wireOut[39]), .ctrl(ctrl[19]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_20(.inData_0(wireIn[40]), .inData_1(wireIn[41]), .outData_0(wireOut[40]), .outData_1(wireOut[41]), .ctrl(ctrl[20]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_21(.inData_0(wireIn[42]), .inData_1(wireIn[43]), .outData_0(wireOut[42]), .outData_1(wireOut[43]), .ctrl(ctrl[21]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_22(.inData_0(wireIn[44]), .inData_1(wireIn[45]), .outData_0(wireOut[44]), .outData_1(wireOut[45]), .ctrl(ctrl[22]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_23(.inData_0(wireIn[46]), .inData_1(wireIn[47]), .outData_0(wireOut[46]), .outData_1(wireOut[47]), .ctrl(ctrl[23]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_24(.inData_0(wireIn[48]), .inData_1(wireIn[49]), .outData_0(wireOut[48]), .outData_1(wireOut[49]), .ctrl(ctrl[24]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_25(.inData_0(wireIn[50]), .inData_1(wireIn[51]), .outData_0(wireOut[50]), .outData_1(wireOut[51]), .ctrl(ctrl[25]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_26(.inData_0(wireIn[52]), .inData_1(wireIn[53]), .outData_0(wireOut[52]), .outData_1(wireOut[53]), .ctrl(ctrl[26]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_27(.inData_0(wireIn[54]), .inData_1(wireIn[55]), .outData_0(wireOut[54]), .outData_1(wireOut[55]), .ctrl(ctrl[27]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_28(.inData_0(wireIn[56]), .inData_1(wireIn[57]), .outData_0(wireOut[56]), .outData_1(wireOut[57]), .ctrl(ctrl[28]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_29(.inData_0(wireIn[58]), .inData_1(wireIn[59]), .outData_0(wireOut[58]), .outData_1(wireOut[59]), .ctrl(ctrl[29]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_30(.inData_0(wireIn[60]), .inData_1(wireIn[61]), .outData_0(wireOut[60]), .outData_1(wireOut[61]), .ctrl(ctrl[30]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_31(.inData_0(wireIn[62]), .inData_1(wireIn[63]), .outData_0(wireOut[62]), .outData_1(wireOut[63]), .ctrl(ctrl[31]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_32(.inData_0(wireIn[64]), .inData_1(wireIn[65]), .outData_0(wireOut[64]), .outData_1(wireOut[65]), .ctrl(ctrl[32]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_33(.inData_0(wireIn[66]), .inData_1(wireIn[67]), .outData_0(wireOut[66]), .outData_1(wireOut[67]), .ctrl(ctrl[33]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_34(.inData_0(wireIn[68]), .inData_1(wireIn[69]), .outData_0(wireOut[68]), .outData_1(wireOut[69]), .ctrl(ctrl[34]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_35(.inData_0(wireIn[70]), .inData_1(wireIn[71]), .outData_0(wireOut[70]), .outData_1(wireOut[71]), .ctrl(ctrl[35]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_36(.inData_0(wireIn[72]), .inData_1(wireIn[73]), .outData_0(wireOut[72]), .outData_1(wireOut[73]), .ctrl(ctrl[36]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_37(.inData_0(wireIn[74]), .inData_1(wireIn[75]), .outData_0(wireOut[74]), .outData_1(wireOut[75]), .ctrl(ctrl[37]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_38(.inData_0(wireIn[76]), .inData_1(wireIn[77]), .outData_0(wireOut[76]), .outData_1(wireOut[77]), .ctrl(ctrl[38]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_39(.inData_0(wireIn[78]), .inData_1(wireIn[79]), .outData_0(wireOut[78]), .outData_1(wireOut[79]), .ctrl(ctrl[39]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_40(.inData_0(wireIn[80]), .inData_1(wireIn[81]), .outData_0(wireOut[80]), .outData_1(wireOut[81]), .ctrl(ctrl[40]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_41(.inData_0(wireIn[82]), .inData_1(wireIn[83]), .outData_0(wireOut[82]), .outData_1(wireOut[83]), .ctrl(ctrl[41]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_42(.inData_0(wireIn[84]), .inData_1(wireIn[85]), .outData_0(wireOut[84]), .outData_1(wireOut[85]), .ctrl(ctrl[42]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_43(.inData_0(wireIn[86]), .inData_1(wireIn[87]), .outData_0(wireOut[86]), .outData_1(wireOut[87]), .ctrl(ctrl[43]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_44(.inData_0(wireIn[88]), .inData_1(wireIn[89]), .outData_0(wireOut[88]), .outData_1(wireOut[89]), .ctrl(ctrl[44]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_45(.inData_0(wireIn[90]), .inData_1(wireIn[91]), .outData_0(wireOut[90]), .outData_1(wireOut[91]), .ctrl(ctrl[45]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_46(.inData_0(wireIn[92]), .inData_1(wireIn[93]), .outData_0(wireOut[92]), .outData_1(wireOut[93]), .ctrl(ctrl[46]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_47(.inData_0(wireIn[94]), .inData_1(wireIn[95]), .outData_0(wireOut[94]), .outData_1(wireOut[95]), .ctrl(ctrl[47]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_48(.inData_0(wireIn[96]), .inData_1(wireIn[97]), .outData_0(wireOut[96]), .outData_1(wireOut[97]), .ctrl(ctrl[48]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_49(.inData_0(wireIn[98]), .inData_1(wireIn[99]), .outData_0(wireOut[98]), .outData_1(wireOut[99]), .ctrl(ctrl[49]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_50(.inData_0(wireIn[100]), .inData_1(wireIn[101]), .outData_0(wireOut[100]), .outData_1(wireOut[101]), .ctrl(ctrl[50]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_51(.inData_0(wireIn[102]), .inData_1(wireIn[103]), .outData_0(wireOut[102]), .outData_1(wireOut[103]), .ctrl(ctrl[51]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_52(.inData_0(wireIn[104]), .inData_1(wireIn[105]), .outData_0(wireOut[104]), .outData_1(wireOut[105]), .ctrl(ctrl[52]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_53(.inData_0(wireIn[106]), .inData_1(wireIn[107]), .outData_0(wireOut[106]), .outData_1(wireOut[107]), .ctrl(ctrl[53]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_54(.inData_0(wireIn[108]), .inData_1(wireIn[109]), .outData_0(wireOut[108]), .outData_1(wireOut[109]), .ctrl(ctrl[54]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_55(.inData_0(wireIn[110]), .inData_1(wireIn[111]), .outData_0(wireOut[110]), .outData_1(wireOut[111]), .ctrl(ctrl[55]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_56(.inData_0(wireIn[112]), .inData_1(wireIn[113]), .outData_0(wireOut[112]), .outData_1(wireOut[113]), .ctrl(ctrl[56]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_57(.inData_0(wireIn[114]), .inData_1(wireIn[115]), .outData_0(wireOut[114]), .outData_1(wireOut[115]), .ctrl(ctrl[57]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_58(.inData_0(wireIn[116]), .inData_1(wireIn[117]), .outData_0(wireOut[116]), .outData_1(wireOut[117]), .ctrl(ctrl[58]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_59(.inData_0(wireIn[118]), .inData_1(wireIn[119]), .outData_0(wireOut[118]), .outData_1(wireOut[119]), .ctrl(ctrl[59]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_60(.inData_0(wireIn[120]), .inData_1(wireIn[121]), .outData_0(wireOut[120]), .outData_1(wireOut[121]), .ctrl(ctrl[60]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_61(.inData_0(wireIn[122]), .inData_1(wireIn[123]), .outData_0(wireOut[122]), .outData_1(wireOut[123]), .ctrl(ctrl[61]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_62(.inData_0(wireIn[124]), .inData_1(wireIn[125]), .outData_0(wireOut[124]), .outData_1(wireOut[125]), .ctrl(ctrl[62]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_63(.inData_0(wireIn[126]), .inData_1(wireIn[127]), .outData_0(wireOut[126]), .outData_1(wireOut[127]), .ctrl(ctrl[63]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_64(.inData_0(wireIn[128]), .inData_1(wireIn[129]), .outData_0(wireOut[128]), .outData_1(wireOut[129]), .ctrl(ctrl[64]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_65(.inData_0(wireIn[130]), .inData_1(wireIn[131]), .outData_0(wireOut[130]), .outData_1(wireOut[131]), .ctrl(ctrl[65]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_66(.inData_0(wireIn[132]), .inData_1(wireIn[133]), .outData_0(wireOut[132]), .outData_1(wireOut[133]), .ctrl(ctrl[66]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_67(.inData_0(wireIn[134]), .inData_1(wireIn[135]), .outData_0(wireOut[134]), .outData_1(wireOut[135]), .ctrl(ctrl[67]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_68(.inData_0(wireIn[136]), .inData_1(wireIn[137]), .outData_0(wireOut[136]), .outData_1(wireOut[137]), .ctrl(ctrl[68]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_69(.inData_0(wireIn[138]), .inData_1(wireIn[139]), .outData_0(wireOut[138]), .outData_1(wireOut[139]), .ctrl(ctrl[69]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_70(.inData_0(wireIn[140]), .inData_1(wireIn[141]), .outData_0(wireOut[140]), .outData_1(wireOut[141]), .ctrl(ctrl[70]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_71(.inData_0(wireIn[142]), .inData_1(wireIn[143]), .outData_0(wireOut[142]), .outData_1(wireOut[143]), .ctrl(ctrl[71]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_72(.inData_0(wireIn[144]), .inData_1(wireIn[145]), .outData_0(wireOut[144]), .outData_1(wireOut[145]), .ctrl(ctrl[72]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_73(.inData_0(wireIn[146]), .inData_1(wireIn[147]), .outData_0(wireOut[146]), .outData_1(wireOut[147]), .ctrl(ctrl[73]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_74(.inData_0(wireIn[148]), .inData_1(wireIn[149]), .outData_0(wireOut[148]), .outData_1(wireOut[149]), .ctrl(ctrl[74]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_75(.inData_0(wireIn[150]), .inData_1(wireIn[151]), .outData_0(wireOut[150]), .outData_1(wireOut[151]), .ctrl(ctrl[75]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_76(.inData_0(wireIn[152]), .inData_1(wireIn[153]), .outData_0(wireOut[152]), .outData_1(wireOut[153]), .ctrl(ctrl[76]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_77(.inData_0(wireIn[154]), .inData_1(wireIn[155]), .outData_0(wireOut[154]), .outData_1(wireOut[155]), .ctrl(ctrl[77]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_78(.inData_0(wireIn[156]), .inData_1(wireIn[157]), .outData_0(wireOut[156]), .outData_1(wireOut[157]), .ctrl(ctrl[78]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_79(.inData_0(wireIn[158]), .inData_1(wireIn[159]), .outData_0(wireOut[158]), .outData_1(wireOut[159]), .ctrl(ctrl[79]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_80(.inData_0(wireIn[160]), .inData_1(wireIn[161]), .outData_0(wireOut[160]), .outData_1(wireOut[161]), .ctrl(ctrl[80]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_81(.inData_0(wireIn[162]), .inData_1(wireIn[163]), .outData_0(wireOut[162]), .outData_1(wireOut[163]), .ctrl(ctrl[81]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_82(.inData_0(wireIn[164]), .inData_1(wireIn[165]), .outData_0(wireOut[164]), .outData_1(wireOut[165]), .ctrl(ctrl[82]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_83(.inData_0(wireIn[166]), .inData_1(wireIn[167]), .outData_0(wireOut[166]), .outData_1(wireOut[167]), .ctrl(ctrl[83]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_84(.inData_0(wireIn[168]), .inData_1(wireIn[169]), .outData_0(wireOut[168]), .outData_1(wireOut[169]), .ctrl(ctrl[84]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_85(.inData_0(wireIn[170]), .inData_1(wireIn[171]), .outData_0(wireOut[170]), .outData_1(wireOut[171]), .ctrl(ctrl[85]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_86(.inData_0(wireIn[172]), .inData_1(wireIn[173]), .outData_0(wireOut[172]), .outData_1(wireOut[173]), .ctrl(ctrl[86]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_87(.inData_0(wireIn[174]), .inData_1(wireIn[175]), .outData_0(wireOut[174]), .outData_1(wireOut[175]), .ctrl(ctrl[87]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_88(.inData_0(wireIn[176]), .inData_1(wireIn[177]), .outData_0(wireOut[176]), .outData_1(wireOut[177]), .ctrl(ctrl[88]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_89(.inData_0(wireIn[178]), .inData_1(wireIn[179]), .outData_0(wireOut[178]), .outData_1(wireOut[179]), .ctrl(ctrl[89]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_90(.inData_0(wireIn[180]), .inData_1(wireIn[181]), .outData_0(wireOut[180]), .outData_1(wireOut[181]), .ctrl(ctrl[90]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_91(.inData_0(wireIn[182]), .inData_1(wireIn[183]), .outData_0(wireOut[182]), .outData_1(wireOut[183]), .ctrl(ctrl[91]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_92(.inData_0(wireIn[184]), .inData_1(wireIn[185]), .outData_0(wireOut[184]), .outData_1(wireOut[185]), .ctrl(ctrl[92]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_93(.inData_0(wireIn[186]), .inData_1(wireIn[187]), .outData_0(wireOut[186]), .outData_1(wireOut[187]), .ctrl(ctrl[93]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_94(.inData_0(wireIn[188]), .inData_1(wireIn[189]), .outData_0(wireOut[188]), .outData_1(wireOut[189]), .ctrl(ctrl[94]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_95(.inData_0(wireIn[190]), .inData_1(wireIn[191]), .outData_0(wireOut[190]), .outData_1(wireOut[191]), .ctrl(ctrl[95]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_96(.inData_0(wireIn[192]), .inData_1(wireIn[193]), .outData_0(wireOut[192]), .outData_1(wireOut[193]), .ctrl(ctrl[96]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_97(.inData_0(wireIn[194]), .inData_1(wireIn[195]), .outData_0(wireOut[194]), .outData_1(wireOut[195]), .ctrl(ctrl[97]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_98(.inData_0(wireIn[196]), .inData_1(wireIn[197]), .outData_0(wireOut[196]), .outData_1(wireOut[197]), .ctrl(ctrl[98]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_99(.inData_0(wireIn[198]), .inData_1(wireIn[199]), .outData_0(wireOut[198]), .outData_1(wireOut[199]), .ctrl(ctrl[99]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_100(.inData_0(wireIn[200]), .inData_1(wireIn[201]), .outData_0(wireOut[200]), .outData_1(wireOut[201]), .ctrl(ctrl[100]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_101(.inData_0(wireIn[202]), .inData_1(wireIn[203]), .outData_0(wireOut[202]), .outData_1(wireOut[203]), .ctrl(ctrl[101]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_102(.inData_0(wireIn[204]), .inData_1(wireIn[205]), .outData_0(wireOut[204]), .outData_1(wireOut[205]), .ctrl(ctrl[102]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_103(.inData_0(wireIn[206]), .inData_1(wireIn[207]), .outData_0(wireOut[206]), .outData_1(wireOut[207]), .ctrl(ctrl[103]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_104(.inData_0(wireIn[208]), .inData_1(wireIn[209]), .outData_0(wireOut[208]), .outData_1(wireOut[209]), .ctrl(ctrl[104]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_105(.inData_0(wireIn[210]), .inData_1(wireIn[211]), .outData_0(wireOut[210]), .outData_1(wireOut[211]), .ctrl(ctrl[105]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_106(.inData_0(wireIn[212]), .inData_1(wireIn[213]), .outData_0(wireOut[212]), .outData_1(wireOut[213]), .ctrl(ctrl[106]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_107(.inData_0(wireIn[214]), .inData_1(wireIn[215]), .outData_0(wireOut[214]), .outData_1(wireOut[215]), .ctrl(ctrl[107]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_108(.inData_0(wireIn[216]), .inData_1(wireIn[217]), .outData_0(wireOut[216]), .outData_1(wireOut[217]), .ctrl(ctrl[108]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_109(.inData_0(wireIn[218]), .inData_1(wireIn[219]), .outData_0(wireOut[218]), .outData_1(wireOut[219]), .ctrl(ctrl[109]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_110(.inData_0(wireIn[220]), .inData_1(wireIn[221]), .outData_0(wireOut[220]), .outData_1(wireOut[221]), .ctrl(ctrl[110]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_111(.inData_0(wireIn[222]), .inData_1(wireIn[223]), .outData_0(wireOut[222]), .outData_1(wireOut[223]), .ctrl(ctrl[111]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_112(.inData_0(wireIn[224]), .inData_1(wireIn[225]), .outData_0(wireOut[224]), .outData_1(wireOut[225]), .ctrl(ctrl[112]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_113(.inData_0(wireIn[226]), .inData_1(wireIn[227]), .outData_0(wireOut[226]), .outData_1(wireOut[227]), .ctrl(ctrl[113]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_114(.inData_0(wireIn[228]), .inData_1(wireIn[229]), .outData_0(wireOut[228]), .outData_1(wireOut[229]), .ctrl(ctrl[114]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_115(.inData_0(wireIn[230]), .inData_1(wireIn[231]), .outData_0(wireOut[230]), .outData_1(wireOut[231]), .ctrl(ctrl[115]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_116(.inData_0(wireIn[232]), .inData_1(wireIn[233]), .outData_0(wireOut[232]), .outData_1(wireOut[233]), .ctrl(ctrl[116]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_117(.inData_0(wireIn[234]), .inData_1(wireIn[235]), .outData_0(wireOut[234]), .outData_1(wireOut[235]), .ctrl(ctrl[117]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_118(.inData_0(wireIn[236]), .inData_1(wireIn[237]), .outData_0(wireOut[236]), .outData_1(wireOut[237]), .ctrl(ctrl[118]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_119(.inData_0(wireIn[238]), .inData_1(wireIn[239]), .outData_0(wireOut[238]), .outData_1(wireOut[239]), .ctrl(ctrl[119]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_120(.inData_0(wireIn[240]), .inData_1(wireIn[241]), .outData_0(wireOut[240]), .outData_1(wireOut[241]), .ctrl(ctrl[120]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_121(.inData_0(wireIn[242]), .inData_1(wireIn[243]), .outData_0(wireOut[242]), .outData_1(wireOut[243]), .ctrl(ctrl[121]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_122(.inData_0(wireIn[244]), .inData_1(wireIn[245]), .outData_0(wireOut[244]), .outData_1(wireOut[245]), .ctrl(ctrl[122]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_123(.inData_0(wireIn[246]), .inData_1(wireIn[247]), .outData_0(wireOut[246]), .outData_1(wireOut[247]), .ctrl(ctrl[123]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_124(.inData_0(wireIn[248]), .inData_1(wireIn[249]), .outData_0(wireOut[248]), .outData_1(wireOut[249]), .ctrl(ctrl[124]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_125(.inData_0(wireIn[250]), .inData_1(wireIn[251]), .outData_0(wireOut[250]), .outData_1(wireOut[251]), .ctrl(ctrl[125]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_126(.inData_0(wireIn[252]), .inData_1(wireIn[253]), .outData_0(wireOut[252]), .outData_1(wireOut[253]), .ctrl(ctrl[126]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_127(.inData_0(wireIn[254]), .inData_1(wireIn[255]), .outData_0(wireOut[254]), .outData_1(wireOut[255]), .ctrl(ctrl[127]), .clk(clk), .rst(rst));
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module wireCon_dp256_st3_L(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  assign wireOut[0] = wireIn[0];    
  assign wireOut[1] = wireIn[2];    
  assign wireOut[2] = wireIn[4];    
  assign wireOut[3] = wireIn[6];    
  assign wireOut[4] = wireIn[8];    
  assign wireOut[5] = wireIn[10];    
  assign wireOut[6] = wireIn[12];    
  assign wireOut[7] = wireIn[14];    
  assign wireOut[8] = wireIn[16];    
  assign wireOut[9] = wireIn[18];    
  assign wireOut[10] = wireIn[20];    
  assign wireOut[11] = wireIn[22];    
  assign wireOut[12] = wireIn[24];    
  assign wireOut[13] = wireIn[26];    
  assign wireOut[14] = wireIn[28];    
  assign wireOut[15] = wireIn[30];    
  assign wireOut[16] = wireIn[1];    
  assign wireOut[17] = wireIn[3];    
  assign wireOut[18] = wireIn[5];    
  assign wireOut[19] = wireIn[7];    
  assign wireOut[20] = wireIn[9];    
  assign wireOut[21] = wireIn[11];    
  assign wireOut[22] = wireIn[13];    
  assign wireOut[23] = wireIn[15];    
  assign wireOut[24] = wireIn[17];    
  assign wireOut[25] = wireIn[19];    
  assign wireOut[26] = wireIn[21];    
  assign wireOut[27] = wireIn[23];    
  assign wireOut[28] = wireIn[25];    
  assign wireOut[29] = wireIn[27];    
  assign wireOut[30] = wireIn[29];    
  assign wireOut[31] = wireIn[31];    
  assign wireOut[32] = wireIn[32];    
  assign wireOut[33] = wireIn[34];    
  assign wireOut[34] = wireIn[36];    
  assign wireOut[35] = wireIn[38];    
  assign wireOut[36] = wireIn[40];    
  assign wireOut[37] = wireIn[42];    
  assign wireOut[38] = wireIn[44];    
  assign wireOut[39] = wireIn[46];    
  assign wireOut[40] = wireIn[48];    
  assign wireOut[41] = wireIn[50];    
  assign wireOut[42] = wireIn[52];    
  assign wireOut[43] = wireIn[54];    
  assign wireOut[44] = wireIn[56];    
  assign wireOut[45] = wireIn[58];    
  assign wireOut[46] = wireIn[60];    
  assign wireOut[47] = wireIn[62];    
  assign wireOut[48] = wireIn[33];    
  assign wireOut[49] = wireIn[35];    
  assign wireOut[50] = wireIn[37];    
  assign wireOut[51] = wireIn[39];    
  assign wireOut[52] = wireIn[41];    
  assign wireOut[53] = wireIn[43];    
  assign wireOut[54] = wireIn[45];    
  assign wireOut[55] = wireIn[47];    
  assign wireOut[56] = wireIn[49];    
  assign wireOut[57] = wireIn[51];    
  assign wireOut[58] = wireIn[53];    
  assign wireOut[59] = wireIn[55];    
  assign wireOut[60] = wireIn[57];    
  assign wireOut[61] = wireIn[59];    
  assign wireOut[62] = wireIn[61];    
  assign wireOut[63] = wireIn[63];    
  assign wireOut[64] = wireIn[64];    
  assign wireOut[65] = wireIn[66];    
  assign wireOut[66] = wireIn[68];    
  assign wireOut[67] = wireIn[70];    
  assign wireOut[68] = wireIn[72];    
  assign wireOut[69] = wireIn[74];    
  assign wireOut[70] = wireIn[76];    
  assign wireOut[71] = wireIn[78];    
  assign wireOut[72] = wireIn[80];    
  assign wireOut[73] = wireIn[82];    
  assign wireOut[74] = wireIn[84];    
  assign wireOut[75] = wireIn[86];    
  assign wireOut[76] = wireIn[88];    
  assign wireOut[77] = wireIn[90];    
  assign wireOut[78] = wireIn[92];    
  assign wireOut[79] = wireIn[94];    
  assign wireOut[80] = wireIn[65];    
  assign wireOut[81] = wireIn[67];    
  assign wireOut[82] = wireIn[69];    
  assign wireOut[83] = wireIn[71];    
  assign wireOut[84] = wireIn[73];    
  assign wireOut[85] = wireIn[75];    
  assign wireOut[86] = wireIn[77];    
  assign wireOut[87] = wireIn[79];    
  assign wireOut[88] = wireIn[81];    
  assign wireOut[89] = wireIn[83];    
  assign wireOut[90] = wireIn[85];    
  assign wireOut[91] = wireIn[87];    
  assign wireOut[92] = wireIn[89];    
  assign wireOut[93] = wireIn[91];    
  assign wireOut[94] = wireIn[93];    
  assign wireOut[95] = wireIn[95];    
  assign wireOut[96] = wireIn[96];    
  assign wireOut[97] = wireIn[98];    
  assign wireOut[98] = wireIn[100];    
  assign wireOut[99] = wireIn[102];    
  assign wireOut[100] = wireIn[104];    
  assign wireOut[101] = wireIn[106];    
  assign wireOut[102] = wireIn[108];    
  assign wireOut[103] = wireIn[110];    
  assign wireOut[104] = wireIn[112];    
  assign wireOut[105] = wireIn[114];    
  assign wireOut[106] = wireIn[116];    
  assign wireOut[107] = wireIn[118];    
  assign wireOut[108] = wireIn[120];    
  assign wireOut[109] = wireIn[122];    
  assign wireOut[110] = wireIn[124];    
  assign wireOut[111] = wireIn[126];    
  assign wireOut[112] = wireIn[97];    
  assign wireOut[113] = wireIn[99];    
  assign wireOut[114] = wireIn[101];    
  assign wireOut[115] = wireIn[103];    
  assign wireOut[116] = wireIn[105];    
  assign wireOut[117] = wireIn[107];    
  assign wireOut[118] = wireIn[109];    
  assign wireOut[119] = wireIn[111];    
  assign wireOut[120] = wireIn[113];    
  assign wireOut[121] = wireIn[115];    
  assign wireOut[122] = wireIn[117];    
  assign wireOut[123] = wireIn[119];    
  assign wireOut[124] = wireIn[121];    
  assign wireOut[125] = wireIn[123];    
  assign wireOut[126] = wireIn[125];    
  assign wireOut[127] = wireIn[127];    
  assign wireOut[128] = wireIn[128];    
  assign wireOut[129] = wireIn[130];    
  assign wireOut[130] = wireIn[132];    
  assign wireOut[131] = wireIn[134];    
  assign wireOut[132] = wireIn[136];    
  assign wireOut[133] = wireIn[138];    
  assign wireOut[134] = wireIn[140];    
  assign wireOut[135] = wireIn[142];    
  assign wireOut[136] = wireIn[144];    
  assign wireOut[137] = wireIn[146];    
  assign wireOut[138] = wireIn[148];    
  assign wireOut[139] = wireIn[150];    
  assign wireOut[140] = wireIn[152];    
  assign wireOut[141] = wireIn[154];    
  assign wireOut[142] = wireIn[156];    
  assign wireOut[143] = wireIn[158];    
  assign wireOut[144] = wireIn[129];    
  assign wireOut[145] = wireIn[131];    
  assign wireOut[146] = wireIn[133];    
  assign wireOut[147] = wireIn[135];    
  assign wireOut[148] = wireIn[137];    
  assign wireOut[149] = wireIn[139];    
  assign wireOut[150] = wireIn[141];    
  assign wireOut[151] = wireIn[143];    
  assign wireOut[152] = wireIn[145];    
  assign wireOut[153] = wireIn[147];    
  assign wireOut[154] = wireIn[149];    
  assign wireOut[155] = wireIn[151];    
  assign wireOut[156] = wireIn[153];    
  assign wireOut[157] = wireIn[155];    
  assign wireOut[158] = wireIn[157];    
  assign wireOut[159] = wireIn[159];    
  assign wireOut[160] = wireIn[160];    
  assign wireOut[161] = wireIn[162];    
  assign wireOut[162] = wireIn[164];    
  assign wireOut[163] = wireIn[166];    
  assign wireOut[164] = wireIn[168];    
  assign wireOut[165] = wireIn[170];    
  assign wireOut[166] = wireIn[172];    
  assign wireOut[167] = wireIn[174];    
  assign wireOut[168] = wireIn[176];    
  assign wireOut[169] = wireIn[178];    
  assign wireOut[170] = wireIn[180];    
  assign wireOut[171] = wireIn[182];    
  assign wireOut[172] = wireIn[184];    
  assign wireOut[173] = wireIn[186];    
  assign wireOut[174] = wireIn[188];    
  assign wireOut[175] = wireIn[190];    
  assign wireOut[176] = wireIn[161];    
  assign wireOut[177] = wireIn[163];    
  assign wireOut[178] = wireIn[165];    
  assign wireOut[179] = wireIn[167];    
  assign wireOut[180] = wireIn[169];    
  assign wireOut[181] = wireIn[171];    
  assign wireOut[182] = wireIn[173];    
  assign wireOut[183] = wireIn[175];    
  assign wireOut[184] = wireIn[177];    
  assign wireOut[185] = wireIn[179];    
  assign wireOut[186] = wireIn[181];    
  assign wireOut[187] = wireIn[183];    
  assign wireOut[188] = wireIn[185];    
  assign wireOut[189] = wireIn[187];    
  assign wireOut[190] = wireIn[189];    
  assign wireOut[191] = wireIn[191];    
  assign wireOut[192] = wireIn[192];    
  assign wireOut[193] = wireIn[194];    
  assign wireOut[194] = wireIn[196];    
  assign wireOut[195] = wireIn[198];    
  assign wireOut[196] = wireIn[200];    
  assign wireOut[197] = wireIn[202];    
  assign wireOut[198] = wireIn[204];    
  assign wireOut[199] = wireIn[206];    
  assign wireOut[200] = wireIn[208];    
  assign wireOut[201] = wireIn[210];    
  assign wireOut[202] = wireIn[212];    
  assign wireOut[203] = wireIn[214];    
  assign wireOut[204] = wireIn[216];    
  assign wireOut[205] = wireIn[218];    
  assign wireOut[206] = wireIn[220];    
  assign wireOut[207] = wireIn[222];    
  assign wireOut[208] = wireIn[193];    
  assign wireOut[209] = wireIn[195];    
  assign wireOut[210] = wireIn[197];    
  assign wireOut[211] = wireIn[199];    
  assign wireOut[212] = wireIn[201];    
  assign wireOut[213] = wireIn[203];    
  assign wireOut[214] = wireIn[205];    
  assign wireOut[215] = wireIn[207];    
  assign wireOut[216] = wireIn[209];    
  assign wireOut[217] = wireIn[211];    
  assign wireOut[218] = wireIn[213];    
  assign wireOut[219] = wireIn[215];    
  assign wireOut[220] = wireIn[217];    
  assign wireOut[221] = wireIn[219];    
  assign wireOut[222] = wireIn[221];    
  assign wireOut[223] = wireIn[223];    
  assign wireOut[224] = wireIn[224];    
  assign wireOut[225] = wireIn[226];    
  assign wireOut[226] = wireIn[228];    
  assign wireOut[227] = wireIn[230];    
  assign wireOut[228] = wireIn[232];    
  assign wireOut[229] = wireIn[234];    
  assign wireOut[230] = wireIn[236];    
  assign wireOut[231] = wireIn[238];    
  assign wireOut[232] = wireIn[240];    
  assign wireOut[233] = wireIn[242];    
  assign wireOut[234] = wireIn[244];    
  assign wireOut[235] = wireIn[246];    
  assign wireOut[236] = wireIn[248];    
  assign wireOut[237] = wireIn[250];    
  assign wireOut[238] = wireIn[252];    
  assign wireOut[239] = wireIn[254];    
  assign wireOut[240] = wireIn[225];    
  assign wireOut[241] = wireIn[227];    
  assign wireOut[242] = wireIn[229];    
  assign wireOut[243] = wireIn[231];    
  assign wireOut[244] = wireIn[233];    
  assign wireOut[245] = wireIn[235];    
  assign wireOut[246] = wireIn[237];    
  assign wireOut[247] = wireIn[239];    
  assign wireOut[248] = wireIn[241];    
  assign wireOut[249] = wireIn[243];    
  assign wireOut[250] = wireIn[245];    
  assign wireOut[251] = wireIn[247];    
  assign wireOut[252] = wireIn[249];    
  assign wireOut[253] = wireIn[251];    
  assign wireOut[254] = wireIn[253];    
  assign wireOut[255] = wireIn[255];    
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module switches_stage_st4_0_L(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
ctrl,                            
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;                   
  input [128-1:0] ctrl;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  switch_2_2 switch_inst_0(.inData_0(wireIn[0]), .inData_1(wireIn[1]), .outData_0(wireOut[0]), .outData_1(wireOut[1]), .ctrl(ctrl[0]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_1(.inData_0(wireIn[2]), .inData_1(wireIn[3]), .outData_0(wireOut[2]), .outData_1(wireOut[3]), .ctrl(ctrl[1]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_2(.inData_0(wireIn[4]), .inData_1(wireIn[5]), .outData_0(wireOut[4]), .outData_1(wireOut[5]), .ctrl(ctrl[2]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_3(.inData_0(wireIn[6]), .inData_1(wireIn[7]), .outData_0(wireOut[6]), .outData_1(wireOut[7]), .ctrl(ctrl[3]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_4(.inData_0(wireIn[8]), .inData_1(wireIn[9]), .outData_0(wireOut[8]), .outData_1(wireOut[9]), .ctrl(ctrl[4]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_5(.inData_0(wireIn[10]), .inData_1(wireIn[11]), .outData_0(wireOut[10]), .outData_1(wireOut[11]), .ctrl(ctrl[5]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_6(.inData_0(wireIn[12]), .inData_1(wireIn[13]), .outData_0(wireOut[12]), .outData_1(wireOut[13]), .ctrl(ctrl[6]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_7(.inData_0(wireIn[14]), .inData_1(wireIn[15]), .outData_0(wireOut[14]), .outData_1(wireOut[15]), .ctrl(ctrl[7]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_8(.inData_0(wireIn[16]), .inData_1(wireIn[17]), .outData_0(wireOut[16]), .outData_1(wireOut[17]), .ctrl(ctrl[8]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_9(.inData_0(wireIn[18]), .inData_1(wireIn[19]), .outData_0(wireOut[18]), .outData_1(wireOut[19]), .ctrl(ctrl[9]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_10(.inData_0(wireIn[20]), .inData_1(wireIn[21]), .outData_0(wireOut[20]), .outData_1(wireOut[21]), .ctrl(ctrl[10]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_11(.inData_0(wireIn[22]), .inData_1(wireIn[23]), .outData_0(wireOut[22]), .outData_1(wireOut[23]), .ctrl(ctrl[11]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_12(.inData_0(wireIn[24]), .inData_1(wireIn[25]), .outData_0(wireOut[24]), .outData_1(wireOut[25]), .ctrl(ctrl[12]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_13(.inData_0(wireIn[26]), .inData_1(wireIn[27]), .outData_0(wireOut[26]), .outData_1(wireOut[27]), .ctrl(ctrl[13]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_14(.inData_0(wireIn[28]), .inData_1(wireIn[29]), .outData_0(wireOut[28]), .outData_1(wireOut[29]), .ctrl(ctrl[14]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_15(.inData_0(wireIn[30]), .inData_1(wireIn[31]), .outData_0(wireOut[30]), .outData_1(wireOut[31]), .ctrl(ctrl[15]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_16(.inData_0(wireIn[32]), .inData_1(wireIn[33]), .outData_0(wireOut[32]), .outData_1(wireOut[33]), .ctrl(ctrl[16]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_17(.inData_0(wireIn[34]), .inData_1(wireIn[35]), .outData_0(wireOut[34]), .outData_1(wireOut[35]), .ctrl(ctrl[17]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_18(.inData_0(wireIn[36]), .inData_1(wireIn[37]), .outData_0(wireOut[36]), .outData_1(wireOut[37]), .ctrl(ctrl[18]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_19(.inData_0(wireIn[38]), .inData_1(wireIn[39]), .outData_0(wireOut[38]), .outData_1(wireOut[39]), .ctrl(ctrl[19]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_20(.inData_0(wireIn[40]), .inData_1(wireIn[41]), .outData_0(wireOut[40]), .outData_1(wireOut[41]), .ctrl(ctrl[20]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_21(.inData_0(wireIn[42]), .inData_1(wireIn[43]), .outData_0(wireOut[42]), .outData_1(wireOut[43]), .ctrl(ctrl[21]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_22(.inData_0(wireIn[44]), .inData_1(wireIn[45]), .outData_0(wireOut[44]), .outData_1(wireOut[45]), .ctrl(ctrl[22]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_23(.inData_0(wireIn[46]), .inData_1(wireIn[47]), .outData_0(wireOut[46]), .outData_1(wireOut[47]), .ctrl(ctrl[23]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_24(.inData_0(wireIn[48]), .inData_1(wireIn[49]), .outData_0(wireOut[48]), .outData_1(wireOut[49]), .ctrl(ctrl[24]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_25(.inData_0(wireIn[50]), .inData_1(wireIn[51]), .outData_0(wireOut[50]), .outData_1(wireOut[51]), .ctrl(ctrl[25]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_26(.inData_0(wireIn[52]), .inData_1(wireIn[53]), .outData_0(wireOut[52]), .outData_1(wireOut[53]), .ctrl(ctrl[26]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_27(.inData_0(wireIn[54]), .inData_1(wireIn[55]), .outData_0(wireOut[54]), .outData_1(wireOut[55]), .ctrl(ctrl[27]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_28(.inData_0(wireIn[56]), .inData_1(wireIn[57]), .outData_0(wireOut[56]), .outData_1(wireOut[57]), .ctrl(ctrl[28]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_29(.inData_0(wireIn[58]), .inData_1(wireIn[59]), .outData_0(wireOut[58]), .outData_1(wireOut[59]), .ctrl(ctrl[29]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_30(.inData_0(wireIn[60]), .inData_1(wireIn[61]), .outData_0(wireOut[60]), .outData_1(wireOut[61]), .ctrl(ctrl[30]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_31(.inData_0(wireIn[62]), .inData_1(wireIn[63]), .outData_0(wireOut[62]), .outData_1(wireOut[63]), .ctrl(ctrl[31]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_32(.inData_0(wireIn[64]), .inData_1(wireIn[65]), .outData_0(wireOut[64]), .outData_1(wireOut[65]), .ctrl(ctrl[32]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_33(.inData_0(wireIn[66]), .inData_1(wireIn[67]), .outData_0(wireOut[66]), .outData_1(wireOut[67]), .ctrl(ctrl[33]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_34(.inData_0(wireIn[68]), .inData_1(wireIn[69]), .outData_0(wireOut[68]), .outData_1(wireOut[69]), .ctrl(ctrl[34]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_35(.inData_0(wireIn[70]), .inData_1(wireIn[71]), .outData_0(wireOut[70]), .outData_1(wireOut[71]), .ctrl(ctrl[35]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_36(.inData_0(wireIn[72]), .inData_1(wireIn[73]), .outData_0(wireOut[72]), .outData_1(wireOut[73]), .ctrl(ctrl[36]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_37(.inData_0(wireIn[74]), .inData_1(wireIn[75]), .outData_0(wireOut[74]), .outData_1(wireOut[75]), .ctrl(ctrl[37]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_38(.inData_0(wireIn[76]), .inData_1(wireIn[77]), .outData_0(wireOut[76]), .outData_1(wireOut[77]), .ctrl(ctrl[38]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_39(.inData_0(wireIn[78]), .inData_1(wireIn[79]), .outData_0(wireOut[78]), .outData_1(wireOut[79]), .ctrl(ctrl[39]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_40(.inData_0(wireIn[80]), .inData_1(wireIn[81]), .outData_0(wireOut[80]), .outData_1(wireOut[81]), .ctrl(ctrl[40]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_41(.inData_0(wireIn[82]), .inData_1(wireIn[83]), .outData_0(wireOut[82]), .outData_1(wireOut[83]), .ctrl(ctrl[41]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_42(.inData_0(wireIn[84]), .inData_1(wireIn[85]), .outData_0(wireOut[84]), .outData_1(wireOut[85]), .ctrl(ctrl[42]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_43(.inData_0(wireIn[86]), .inData_1(wireIn[87]), .outData_0(wireOut[86]), .outData_1(wireOut[87]), .ctrl(ctrl[43]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_44(.inData_0(wireIn[88]), .inData_1(wireIn[89]), .outData_0(wireOut[88]), .outData_1(wireOut[89]), .ctrl(ctrl[44]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_45(.inData_0(wireIn[90]), .inData_1(wireIn[91]), .outData_0(wireOut[90]), .outData_1(wireOut[91]), .ctrl(ctrl[45]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_46(.inData_0(wireIn[92]), .inData_1(wireIn[93]), .outData_0(wireOut[92]), .outData_1(wireOut[93]), .ctrl(ctrl[46]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_47(.inData_0(wireIn[94]), .inData_1(wireIn[95]), .outData_0(wireOut[94]), .outData_1(wireOut[95]), .ctrl(ctrl[47]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_48(.inData_0(wireIn[96]), .inData_1(wireIn[97]), .outData_0(wireOut[96]), .outData_1(wireOut[97]), .ctrl(ctrl[48]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_49(.inData_0(wireIn[98]), .inData_1(wireIn[99]), .outData_0(wireOut[98]), .outData_1(wireOut[99]), .ctrl(ctrl[49]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_50(.inData_0(wireIn[100]), .inData_1(wireIn[101]), .outData_0(wireOut[100]), .outData_1(wireOut[101]), .ctrl(ctrl[50]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_51(.inData_0(wireIn[102]), .inData_1(wireIn[103]), .outData_0(wireOut[102]), .outData_1(wireOut[103]), .ctrl(ctrl[51]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_52(.inData_0(wireIn[104]), .inData_1(wireIn[105]), .outData_0(wireOut[104]), .outData_1(wireOut[105]), .ctrl(ctrl[52]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_53(.inData_0(wireIn[106]), .inData_1(wireIn[107]), .outData_0(wireOut[106]), .outData_1(wireOut[107]), .ctrl(ctrl[53]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_54(.inData_0(wireIn[108]), .inData_1(wireIn[109]), .outData_0(wireOut[108]), .outData_1(wireOut[109]), .ctrl(ctrl[54]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_55(.inData_0(wireIn[110]), .inData_1(wireIn[111]), .outData_0(wireOut[110]), .outData_1(wireOut[111]), .ctrl(ctrl[55]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_56(.inData_0(wireIn[112]), .inData_1(wireIn[113]), .outData_0(wireOut[112]), .outData_1(wireOut[113]), .ctrl(ctrl[56]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_57(.inData_0(wireIn[114]), .inData_1(wireIn[115]), .outData_0(wireOut[114]), .outData_1(wireOut[115]), .ctrl(ctrl[57]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_58(.inData_0(wireIn[116]), .inData_1(wireIn[117]), .outData_0(wireOut[116]), .outData_1(wireOut[117]), .ctrl(ctrl[58]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_59(.inData_0(wireIn[118]), .inData_1(wireIn[119]), .outData_0(wireOut[118]), .outData_1(wireOut[119]), .ctrl(ctrl[59]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_60(.inData_0(wireIn[120]), .inData_1(wireIn[121]), .outData_0(wireOut[120]), .outData_1(wireOut[121]), .ctrl(ctrl[60]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_61(.inData_0(wireIn[122]), .inData_1(wireIn[123]), .outData_0(wireOut[122]), .outData_1(wireOut[123]), .ctrl(ctrl[61]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_62(.inData_0(wireIn[124]), .inData_1(wireIn[125]), .outData_0(wireOut[124]), .outData_1(wireOut[125]), .ctrl(ctrl[62]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_63(.inData_0(wireIn[126]), .inData_1(wireIn[127]), .outData_0(wireOut[126]), .outData_1(wireOut[127]), .ctrl(ctrl[63]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_64(.inData_0(wireIn[128]), .inData_1(wireIn[129]), .outData_0(wireOut[128]), .outData_1(wireOut[129]), .ctrl(ctrl[64]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_65(.inData_0(wireIn[130]), .inData_1(wireIn[131]), .outData_0(wireOut[130]), .outData_1(wireOut[131]), .ctrl(ctrl[65]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_66(.inData_0(wireIn[132]), .inData_1(wireIn[133]), .outData_0(wireOut[132]), .outData_1(wireOut[133]), .ctrl(ctrl[66]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_67(.inData_0(wireIn[134]), .inData_1(wireIn[135]), .outData_0(wireOut[134]), .outData_1(wireOut[135]), .ctrl(ctrl[67]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_68(.inData_0(wireIn[136]), .inData_1(wireIn[137]), .outData_0(wireOut[136]), .outData_1(wireOut[137]), .ctrl(ctrl[68]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_69(.inData_0(wireIn[138]), .inData_1(wireIn[139]), .outData_0(wireOut[138]), .outData_1(wireOut[139]), .ctrl(ctrl[69]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_70(.inData_0(wireIn[140]), .inData_1(wireIn[141]), .outData_0(wireOut[140]), .outData_1(wireOut[141]), .ctrl(ctrl[70]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_71(.inData_0(wireIn[142]), .inData_1(wireIn[143]), .outData_0(wireOut[142]), .outData_1(wireOut[143]), .ctrl(ctrl[71]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_72(.inData_0(wireIn[144]), .inData_1(wireIn[145]), .outData_0(wireOut[144]), .outData_1(wireOut[145]), .ctrl(ctrl[72]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_73(.inData_0(wireIn[146]), .inData_1(wireIn[147]), .outData_0(wireOut[146]), .outData_1(wireOut[147]), .ctrl(ctrl[73]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_74(.inData_0(wireIn[148]), .inData_1(wireIn[149]), .outData_0(wireOut[148]), .outData_1(wireOut[149]), .ctrl(ctrl[74]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_75(.inData_0(wireIn[150]), .inData_1(wireIn[151]), .outData_0(wireOut[150]), .outData_1(wireOut[151]), .ctrl(ctrl[75]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_76(.inData_0(wireIn[152]), .inData_1(wireIn[153]), .outData_0(wireOut[152]), .outData_1(wireOut[153]), .ctrl(ctrl[76]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_77(.inData_0(wireIn[154]), .inData_1(wireIn[155]), .outData_0(wireOut[154]), .outData_1(wireOut[155]), .ctrl(ctrl[77]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_78(.inData_0(wireIn[156]), .inData_1(wireIn[157]), .outData_0(wireOut[156]), .outData_1(wireOut[157]), .ctrl(ctrl[78]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_79(.inData_0(wireIn[158]), .inData_1(wireIn[159]), .outData_0(wireOut[158]), .outData_1(wireOut[159]), .ctrl(ctrl[79]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_80(.inData_0(wireIn[160]), .inData_1(wireIn[161]), .outData_0(wireOut[160]), .outData_1(wireOut[161]), .ctrl(ctrl[80]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_81(.inData_0(wireIn[162]), .inData_1(wireIn[163]), .outData_0(wireOut[162]), .outData_1(wireOut[163]), .ctrl(ctrl[81]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_82(.inData_0(wireIn[164]), .inData_1(wireIn[165]), .outData_0(wireOut[164]), .outData_1(wireOut[165]), .ctrl(ctrl[82]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_83(.inData_0(wireIn[166]), .inData_1(wireIn[167]), .outData_0(wireOut[166]), .outData_1(wireOut[167]), .ctrl(ctrl[83]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_84(.inData_0(wireIn[168]), .inData_1(wireIn[169]), .outData_0(wireOut[168]), .outData_1(wireOut[169]), .ctrl(ctrl[84]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_85(.inData_0(wireIn[170]), .inData_1(wireIn[171]), .outData_0(wireOut[170]), .outData_1(wireOut[171]), .ctrl(ctrl[85]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_86(.inData_0(wireIn[172]), .inData_1(wireIn[173]), .outData_0(wireOut[172]), .outData_1(wireOut[173]), .ctrl(ctrl[86]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_87(.inData_0(wireIn[174]), .inData_1(wireIn[175]), .outData_0(wireOut[174]), .outData_1(wireOut[175]), .ctrl(ctrl[87]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_88(.inData_0(wireIn[176]), .inData_1(wireIn[177]), .outData_0(wireOut[176]), .outData_1(wireOut[177]), .ctrl(ctrl[88]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_89(.inData_0(wireIn[178]), .inData_1(wireIn[179]), .outData_0(wireOut[178]), .outData_1(wireOut[179]), .ctrl(ctrl[89]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_90(.inData_0(wireIn[180]), .inData_1(wireIn[181]), .outData_0(wireOut[180]), .outData_1(wireOut[181]), .ctrl(ctrl[90]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_91(.inData_0(wireIn[182]), .inData_1(wireIn[183]), .outData_0(wireOut[182]), .outData_1(wireOut[183]), .ctrl(ctrl[91]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_92(.inData_0(wireIn[184]), .inData_1(wireIn[185]), .outData_0(wireOut[184]), .outData_1(wireOut[185]), .ctrl(ctrl[92]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_93(.inData_0(wireIn[186]), .inData_1(wireIn[187]), .outData_0(wireOut[186]), .outData_1(wireOut[187]), .ctrl(ctrl[93]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_94(.inData_0(wireIn[188]), .inData_1(wireIn[189]), .outData_0(wireOut[188]), .outData_1(wireOut[189]), .ctrl(ctrl[94]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_95(.inData_0(wireIn[190]), .inData_1(wireIn[191]), .outData_0(wireOut[190]), .outData_1(wireOut[191]), .ctrl(ctrl[95]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_96(.inData_0(wireIn[192]), .inData_1(wireIn[193]), .outData_0(wireOut[192]), .outData_1(wireOut[193]), .ctrl(ctrl[96]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_97(.inData_0(wireIn[194]), .inData_1(wireIn[195]), .outData_0(wireOut[194]), .outData_1(wireOut[195]), .ctrl(ctrl[97]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_98(.inData_0(wireIn[196]), .inData_1(wireIn[197]), .outData_0(wireOut[196]), .outData_1(wireOut[197]), .ctrl(ctrl[98]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_99(.inData_0(wireIn[198]), .inData_1(wireIn[199]), .outData_0(wireOut[198]), .outData_1(wireOut[199]), .ctrl(ctrl[99]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_100(.inData_0(wireIn[200]), .inData_1(wireIn[201]), .outData_0(wireOut[200]), .outData_1(wireOut[201]), .ctrl(ctrl[100]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_101(.inData_0(wireIn[202]), .inData_1(wireIn[203]), .outData_0(wireOut[202]), .outData_1(wireOut[203]), .ctrl(ctrl[101]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_102(.inData_0(wireIn[204]), .inData_1(wireIn[205]), .outData_0(wireOut[204]), .outData_1(wireOut[205]), .ctrl(ctrl[102]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_103(.inData_0(wireIn[206]), .inData_1(wireIn[207]), .outData_0(wireOut[206]), .outData_1(wireOut[207]), .ctrl(ctrl[103]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_104(.inData_0(wireIn[208]), .inData_1(wireIn[209]), .outData_0(wireOut[208]), .outData_1(wireOut[209]), .ctrl(ctrl[104]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_105(.inData_0(wireIn[210]), .inData_1(wireIn[211]), .outData_0(wireOut[210]), .outData_1(wireOut[211]), .ctrl(ctrl[105]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_106(.inData_0(wireIn[212]), .inData_1(wireIn[213]), .outData_0(wireOut[212]), .outData_1(wireOut[213]), .ctrl(ctrl[106]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_107(.inData_0(wireIn[214]), .inData_1(wireIn[215]), .outData_0(wireOut[214]), .outData_1(wireOut[215]), .ctrl(ctrl[107]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_108(.inData_0(wireIn[216]), .inData_1(wireIn[217]), .outData_0(wireOut[216]), .outData_1(wireOut[217]), .ctrl(ctrl[108]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_109(.inData_0(wireIn[218]), .inData_1(wireIn[219]), .outData_0(wireOut[218]), .outData_1(wireOut[219]), .ctrl(ctrl[109]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_110(.inData_0(wireIn[220]), .inData_1(wireIn[221]), .outData_0(wireOut[220]), .outData_1(wireOut[221]), .ctrl(ctrl[110]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_111(.inData_0(wireIn[222]), .inData_1(wireIn[223]), .outData_0(wireOut[222]), .outData_1(wireOut[223]), .ctrl(ctrl[111]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_112(.inData_0(wireIn[224]), .inData_1(wireIn[225]), .outData_0(wireOut[224]), .outData_1(wireOut[225]), .ctrl(ctrl[112]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_113(.inData_0(wireIn[226]), .inData_1(wireIn[227]), .outData_0(wireOut[226]), .outData_1(wireOut[227]), .ctrl(ctrl[113]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_114(.inData_0(wireIn[228]), .inData_1(wireIn[229]), .outData_0(wireOut[228]), .outData_1(wireOut[229]), .ctrl(ctrl[114]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_115(.inData_0(wireIn[230]), .inData_1(wireIn[231]), .outData_0(wireOut[230]), .outData_1(wireOut[231]), .ctrl(ctrl[115]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_116(.inData_0(wireIn[232]), .inData_1(wireIn[233]), .outData_0(wireOut[232]), .outData_1(wireOut[233]), .ctrl(ctrl[116]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_117(.inData_0(wireIn[234]), .inData_1(wireIn[235]), .outData_0(wireOut[234]), .outData_1(wireOut[235]), .ctrl(ctrl[117]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_118(.inData_0(wireIn[236]), .inData_1(wireIn[237]), .outData_0(wireOut[236]), .outData_1(wireOut[237]), .ctrl(ctrl[118]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_119(.inData_0(wireIn[238]), .inData_1(wireIn[239]), .outData_0(wireOut[238]), .outData_1(wireOut[239]), .ctrl(ctrl[119]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_120(.inData_0(wireIn[240]), .inData_1(wireIn[241]), .outData_0(wireOut[240]), .outData_1(wireOut[241]), .ctrl(ctrl[120]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_121(.inData_0(wireIn[242]), .inData_1(wireIn[243]), .outData_0(wireOut[242]), .outData_1(wireOut[243]), .ctrl(ctrl[121]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_122(.inData_0(wireIn[244]), .inData_1(wireIn[245]), .outData_0(wireOut[244]), .outData_1(wireOut[245]), .ctrl(ctrl[122]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_123(.inData_0(wireIn[246]), .inData_1(wireIn[247]), .outData_0(wireOut[246]), .outData_1(wireOut[247]), .ctrl(ctrl[123]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_124(.inData_0(wireIn[248]), .inData_1(wireIn[249]), .outData_0(wireOut[248]), .outData_1(wireOut[249]), .ctrl(ctrl[124]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_125(.inData_0(wireIn[250]), .inData_1(wireIn[251]), .outData_0(wireOut[250]), .outData_1(wireOut[251]), .ctrl(ctrl[125]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_126(.inData_0(wireIn[252]), .inData_1(wireIn[253]), .outData_0(wireOut[252]), .outData_1(wireOut[253]), .ctrl(ctrl[126]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_127(.inData_0(wireIn[254]), .inData_1(wireIn[255]), .outData_0(wireOut[254]), .outData_1(wireOut[255]), .ctrl(ctrl[127]), .clk(clk), .rst(rst));
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module wireCon_dp256_st4_L(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  assign wireOut[0] = wireIn[0];    
  assign wireOut[1] = wireIn[2];    
  assign wireOut[2] = wireIn[4];    
  assign wireOut[3] = wireIn[6];    
  assign wireOut[4] = wireIn[8];    
  assign wireOut[5] = wireIn[10];    
  assign wireOut[6] = wireIn[12];    
  assign wireOut[7] = wireIn[14];    
  assign wireOut[8] = wireIn[1];    
  assign wireOut[9] = wireIn[3];    
  assign wireOut[10] = wireIn[5];    
  assign wireOut[11] = wireIn[7];    
  assign wireOut[12] = wireIn[9];    
  assign wireOut[13] = wireIn[11];    
  assign wireOut[14] = wireIn[13];    
  assign wireOut[15] = wireIn[15];    
  assign wireOut[16] = wireIn[16];    
  assign wireOut[17] = wireIn[18];    
  assign wireOut[18] = wireIn[20];    
  assign wireOut[19] = wireIn[22];    
  assign wireOut[20] = wireIn[24];    
  assign wireOut[21] = wireIn[26];    
  assign wireOut[22] = wireIn[28];    
  assign wireOut[23] = wireIn[30];    
  assign wireOut[24] = wireIn[17];    
  assign wireOut[25] = wireIn[19];    
  assign wireOut[26] = wireIn[21];    
  assign wireOut[27] = wireIn[23];    
  assign wireOut[28] = wireIn[25];    
  assign wireOut[29] = wireIn[27];    
  assign wireOut[30] = wireIn[29];    
  assign wireOut[31] = wireIn[31];    
  assign wireOut[32] = wireIn[32];    
  assign wireOut[33] = wireIn[34];    
  assign wireOut[34] = wireIn[36];    
  assign wireOut[35] = wireIn[38];    
  assign wireOut[36] = wireIn[40];    
  assign wireOut[37] = wireIn[42];    
  assign wireOut[38] = wireIn[44];    
  assign wireOut[39] = wireIn[46];    
  assign wireOut[40] = wireIn[33];    
  assign wireOut[41] = wireIn[35];    
  assign wireOut[42] = wireIn[37];    
  assign wireOut[43] = wireIn[39];    
  assign wireOut[44] = wireIn[41];    
  assign wireOut[45] = wireIn[43];    
  assign wireOut[46] = wireIn[45];    
  assign wireOut[47] = wireIn[47];    
  assign wireOut[48] = wireIn[48];    
  assign wireOut[49] = wireIn[50];    
  assign wireOut[50] = wireIn[52];    
  assign wireOut[51] = wireIn[54];    
  assign wireOut[52] = wireIn[56];    
  assign wireOut[53] = wireIn[58];    
  assign wireOut[54] = wireIn[60];    
  assign wireOut[55] = wireIn[62];    
  assign wireOut[56] = wireIn[49];    
  assign wireOut[57] = wireIn[51];    
  assign wireOut[58] = wireIn[53];    
  assign wireOut[59] = wireIn[55];    
  assign wireOut[60] = wireIn[57];    
  assign wireOut[61] = wireIn[59];    
  assign wireOut[62] = wireIn[61];    
  assign wireOut[63] = wireIn[63];    
  assign wireOut[64] = wireIn[64];    
  assign wireOut[65] = wireIn[66];    
  assign wireOut[66] = wireIn[68];    
  assign wireOut[67] = wireIn[70];    
  assign wireOut[68] = wireIn[72];    
  assign wireOut[69] = wireIn[74];    
  assign wireOut[70] = wireIn[76];    
  assign wireOut[71] = wireIn[78];    
  assign wireOut[72] = wireIn[65];    
  assign wireOut[73] = wireIn[67];    
  assign wireOut[74] = wireIn[69];    
  assign wireOut[75] = wireIn[71];    
  assign wireOut[76] = wireIn[73];    
  assign wireOut[77] = wireIn[75];    
  assign wireOut[78] = wireIn[77];    
  assign wireOut[79] = wireIn[79];    
  assign wireOut[80] = wireIn[80];    
  assign wireOut[81] = wireIn[82];    
  assign wireOut[82] = wireIn[84];    
  assign wireOut[83] = wireIn[86];    
  assign wireOut[84] = wireIn[88];    
  assign wireOut[85] = wireIn[90];    
  assign wireOut[86] = wireIn[92];    
  assign wireOut[87] = wireIn[94];    
  assign wireOut[88] = wireIn[81];    
  assign wireOut[89] = wireIn[83];    
  assign wireOut[90] = wireIn[85];    
  assign wireOut[91] = wireIn[87];    
  assign wireOut[92] = wireIn[89];    
  assign wireOut[93] = wireIn[91];    
  assign wireOut[94] = wireIn[93];    
  assign wireOut[95] = wireIn[95];    
  assign wireOut[96] = wireIn[96];    
  assign wireOut[97] = wireIn[98];    
  assign wireOut[98] = wireIn[100];    
  assign wireOut[99] = wireIn[102];    
  assign wireOut[100] = wireIn[104];    
  assign wireOut[101] = wireIn[106];    
  assign wireOut[102] = wireIn[108];    
  assign wireOut[103] = wireIn[110];    
  assign wireOut[104] = wireIn[97];    
  assign wireOut[105] = wireIn[99];    
  assign wireOut[106] = wireIn[101];    
  assign wireOut[107] = wireIn[103];    
  assign wireOut[108] = wireIn[105];    
  assign wireOut[109] = wireIn[107];    
  assign wireOut[110] = wireIn[109];    
  assign wireOut[111] = wireIn[111];    
  assign wireOut[112] = wireIn[112];    
  assign wireOut[113] = wireIn[114];    
  assign wireOut[114] = wireIn[116];    
  assign wireOut[115] = wireIn[118];    
  assign wireOut[116] = wireIn[120];    
  assign wireOut[117] = wireIn[122];    
  assign wireOut[118] = wireIn[124];    
  assign wireOut[119] = wireIn[126];    
  assign wireOut[120] = wireIn[113];    
  assign wireOut[121] = wireIn[115];    
  assign wireOut[122] = wireIn[117];    
  assign wireOut[123] = wireIn[119];    
  assign wireOut[124] = wireIn[121];    
  assign wireOut[125] = wireIn[123];    
  assign wireOut[126] = wireIn[125];    
  assign wireOut[127] = wireIn[127];    
  assign wireOut[128] = wireIn[128];    
  assign wireOut[129] = wireIn[130];    
  assign wireOut[130] = wireIn[132];    
  assign wireOut[131] = wireIn[134];    
  assign wireOut[132] = wireIn[136];    
  assign wireOut[133] = wireIn[138];    
  assign wireOut[134] = wireIn[140];    
  assign wireOut[135] = wireIn[142];    
  assign wireOut[136] = wireIn[129];    
  assign wireOut[137] = wireIn[131];    
  assign wireOut[138] = wireIn[133];    
  assign wireOut[139] = wireIn[135];    
  assign wireOut[140] = wireIn[137];    
  assign wireOut[141] = wireIn[139];    
  assign wireOut[142] = wireIn[141];    
  assign wireOut[143] = wireIn[143];    
  assign wireOut[144] = wireIn[144];    
  assign wireOut[145] = wireIn[146];    
  assign wireOut[146] = wireIn[148];    
  assign wireOut[147] = wireIn[150];    
  assign wireOut[148] = wireIn[152];    
  assign wireOut[149] = wireIn[154];    
  assign wireOut[150] = wireIn[156];    
  assign wireOut[151] = wireIn[158];    
  assign wireOut[152] = wireIn[145];    
  assign wireOut[153] = wireIn[147];    
  assign wireOut[154] = wireIn[149];    
  assign wireOut[155] = wireIn[151];    
  assign wireOut[156] = wireIn[153];    
  assign wireOut[157] = wireIn[155];    
  assign wireOut[158] = wireIn[157];    
  assign wireOut[159] = wireIn[159];    
  assign wireOut[160] = wireIn[160];    
  assign wireOut[161] = wireIn[162];    
  assign wireOut[162] = wireIn[164];    
  assign wireOut[163] = wireIn[166];    
  assign wireOut[164] = wireIn[168];    
  assign wireOut[165] = wireIn[170];    
  assign wireOut[166] = wireIn[172];    
  assign wireOut[167] = wireIn[174];    
  assign wireOut[168] = wireIn[161];    
  assign wireOut[169] = wireIn[163];    
  assign wireOut[170] = wireIn[165];    
  assign wireOut[171] = wireIn[167];    
  assign wireOut[172] = wireIn[169];    
  assign wireOut[173] = wireIn[171];    
  assign wireOut[174] = wireIn[173];    
  assign wireOut[175] = wireIn[175];    
  assign wireOut[176] = wireIn[176];    
  assign wireOut[177] = wireIn[178];    
  assign wireOut[178] = wireIn[180];    
  assign wireOut[179] = wireIn[182];    
  assign wireOut[180] = wireIn[184];    
  assign wireOut[181] = wireIn[186];    
  assign wireOut[182] = wireIn[188];    
  assign wireOut[183] = wireIn[190];    
  assign wireOut[184] = wireIn[177];    
  assign wireOut[185] = wireIn[179];    
  assign wireOut[186] = wireIn[181];    
  assign wireOut[187] = wireIn[183];    
  assign wireOut[188] = wireIn[185];    
  assign wireOut[189] = wireIn[187];    
  assign wireOut[190] = wireIn[189];    
  assign wireOut[191] = wireIn[191];    
  assign wireOut[192] = wireIn[192];    
  assign wireOut[193] = wireIn[194];    
  assign wireOut[194] = wireIn[196];    
  assign wireOut[195] = wireIn[198];    
  assign wireOut[196] = wireIn[200];    
  assign wireOut[197] = wireIn[202];    
  assign wireOut[198] = wireIn[204];    
  assign wireOut[199] = wireIn[206];    
  assign wireOut[200] = wireIn[193];    
  assign wireOut[201] = wireIn[195];    
  assign wireOut[202] = wireIn[197];    
  assign wireOut[203] = wireIn[199];    
  assign wireOut[204] = wireIn[201];    
  assign wireOut[205] = wireIn[203];    
  assign wireOut[206] = wireIn[205];    
  assign wireOut[207] = wireIn[207];    
  assign wireOut[208] = wireIn[208];    
  assign wireOut[209] = wireIn[210];    
  assign wireOut[210] = wireIn[212];    
  assign wireOut[211] = wireIn[214];    
  assign wireOut[212] = wireIn[216];    
  assign wireOut[213] = wireIn[218];    
  assign wireOut[214] = wireIn[220];    
  assign wireOut[215] = wireIn[222];    
  assign wireOut[216] = wireIn[209];    
  assign wireOut[217] = wireIn[211];    
  assign wireOut[218] = wireIn[213];    
  assign wireOut[219] = wireIn[215];    
  assign wireOut[220] = wireIn[217];    
  assign wireOut[221] = wireIn[219];    
  assign wireOut[222] = wireIn[221];    
  assign wireOut[223] = wireIn[223];    
  assign wireOut[224] = wireIn[224];    
  assign wireOut[225] = wireIn[226];    
  assign wireOut[226] = wireIn[228];    
  assign wireOut[227] = wireIn[230];    
  assign wireOut[228] = wireIn[232];    
  assign wireOut[229] = wireIn[234];    
  assign wireOut[230] = wireIn[236];    
  assign wireOut[231] = wireIn[238];    
  assign wireOut[232] = wireIn[225];    
  assign wireOut[233] = wireIn[227];    
  assign wireOut[234] = wireIn[229];    
  assign wireOut[235] = wireIn[231];    
  assign wireOut[236] = wireIn[233];    
  assign wireOut[237] = wireIn[235];    
  assign wireOut[238] = wireIn[237];    
  assign wireOut[239] = wireIn[239];    
  assign wireOut[240] = wireIn[240];    
  assign wireOut[241] = wireIn[242];    
  assign wireOut[242] = wireIn[244];    
  assign wireOut[243] = wireIn[246];    
  assign wireOut[244] = wireIn[248];    
  assign wireOut[245] = wireIn[250];    
  assign wireOut[246] = wireIn[252];    
  assign wireOut[247] = wireIn[254];    
  assign wireOut[248] = wireIn[241];    
  assign wireOut[249] = wireIn[243];    
  assign wireOut[250] = wireIn[245];    
  assign wireOut[251] = wireIn[247];    
  assign wireOut[252] = wireIn[249];    
  assign wireOut[253] = wireIn[251];    
  assign wireOut[254] = wireIn[253];    
  assign wireOut[255] = wireIn[255];    
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module switches_stage_st5_0_L(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
ctrl,                            
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;                   
  input [128-1:0] ctrl;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  switch_2_2 switch_inst_0(.inData_0(wireIn[0]), .inData_1(wireIn[1]), .outData_0(wireOut[0]), .outData_1(wireOut[1]), .ctrl(ctrl[0]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_1(.inData_0(wireIn[2]), .inData_1(wireIn[3]), .outData_0(wireOut[2]), .outData_1(wireOut[3]), .ctrl(ctrl[1]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_2(.inData_0(wireIn[4]), .inData_1(wireIn[5]), .outData_0(wireOut[4]), .outData_1(wireOut[5]), .ctrl(ctrl[2]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_3(.inData_0(wireIn[6]), .inData_1(wireIn[7]), .outData_0(wireOut[6]), .outData_1(wireOut[7]), .ctrl(ctrl[3]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_4(.inData_0(wireIn[8]), .inData_1(wireIn[9]), .outData_0(wireOut[8]), .outData_1(wireOut[9]), .ctrl(ctrl[4]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_5(.inData_0(wireIn[10]), .inData_1(wireIn[11]), .outData_0(wireOut[10]), .outData_1(wireOut[11]), .ctrl(ctrl[5]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_6(.inData_0(wireIn[12]), .inData_1(wireIn[13]), .outData_0(wireOut[12]), .outData_1(wireOut[13]), .ctrl(ctrl[6]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_7(.inData_0(wireIn[14]), .inData_1(wireIn[15]), .outData_0(wireOut[14]), .outData_1(wireOut[15]), .ctrl(ctrl[7]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_8(.inData_0(wireIn[16]), .inData_1(wireIn[17]), .outData_0(wireOut[16]), .outData_1(wireOut[17]), .ctrl(ctrl[8]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_9(.inData_0(wireIn[18]), .inData_1(wireIn[19]), .outData_0(wireOut[18]), .outData_1(wireOut[19]), .ctrl(ctrl[9]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_10(.inData_0(wireIn[20]), .inData_1(wireIn[21]), .outData_0(wireOut[20]), .outData_1(wireOut[21]), .ctrl(ctrl[10]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_11(.inData_0(wireIn[22]), .inData_1(wireIn[23]), .outData_0(wireOut[22]), .outData_1(wireOut[23]), .ctrl(ctrl[11]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_12(.inData_0(wireIn[24]), .inData_1(wireIn[25]), .outData_0(wireOut[24]), .outData_1(wireOut[25]), .ctrl(ctrl[12]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_13(.inData_0(wireIn[26]), .inData_1(wireIn[27]), .outData_0(wireOut[26]), .outData_1(wireOut[27]), .ctrl(ctrl[13]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_14(.inData_0(wireIn[28]), .inData_1(wireIn[29]), .outData_0(wireOut[28]), .outData_1(wireOut[29]), .ctrl(ctrl[14]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_15(.inData_0(wireIn[30]), .inData_1(wireIn[31]), .outData_0(wireOut[30]), .outData_1(wireOut[31]), .ctrl(ctrl[15]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_16(.inData_0(wireIn[32]), .inData_1(wireIn[33]), .outData_0(wireOut[32]), .outData_1(wireOut[33]), .ctrl(ctrl[16]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_17(.inData_0(wireIn[34]), .inData_1(wireIn[35]), .outData_0(wireOut[34]), .outData_1(wireOut[35]), .ctrl(ctrl[17]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_18(.inData_0(wireIn[36]), .inData_1(wireIn[37]), .outData_0(wireOut[36]), .outData_1(wireOut[37]), .ctrl(ctrl[18]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_19(.inData_0(wireIn[38]), .inData_1(wireIn[39]), .outData_0(wireOut[38]), .outData_1(wireOut[39]), .ctrl(ctrl[19]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_20(.inData_0(wireIn[40]), .inData_1(wireIn[41]), .outData_0(wireOut[40]), .outData_1(wireOut[41]), .ctrl(ctrl[20]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_21(.inData_0(wireIn[42]), .inData_1(wireIn[43]), .outData_0(wireOut[42]), .outData_1(wireOut[43]), .ctrl(ctrl[21]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_22(.inData_0(wireIn[44]), .inData_1(wireIn[45]), .outData_0(wireOut[44]), .outData_1(wireOut[45]), .ctrl(ctrl[22]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_23(.inData_0(wireIn[46]), .inData_1(wireIn[47]), .outData_0(wireOut[46]), .outData_1(wireOut[47]), .ctrl(ctrl[23]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_24(.inData_0(wireIn[48]), .inData_1(wireIn[49]), .outData_0(wireOut[48]), .outData_1(wireOut[49]), .ctrl(ctrl[24]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_25(.inData_0(wireIn[50]), .inData_1(wireIn[51]), .outData_0(wireOut[50]), .outData_1(wireOut[51]), .ctrl(ctrl[25]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_26(.inData_0(wireIn[52]), .inData_1(wireIn[53]), .outData_0(wireOut[52]), .outData_1(wireOut[53]), .ctrl(ctrl[26]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_27(.inData_0(wireIn[54]), .inData_1(wireIn[55]), .outData_0(wireOut[54]), .outData_1(wireOut[55]), .ctrl(ctrl[27]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_28(.inData_0(wireIn[56]), .inData_1(wireIn[57]), .outData_0(wireOut[56]), .outData_1(wireOut[57]), .ctrl(ctrl[28]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_29(.inData_0(wireIn[58]), .inData_1(wireIn[59]), .outData_0(wireOut[58]), .outData_1(wireOut[59]), .ctrl(ctrl[29]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_30(.inData_0(wireIn[60]), .inData_1(wireIn[61]), .outData_0(wireOut[60]), .outData_1(wireOut[61]), .ctrl(ctrl[30]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_31(.inData_0(wireIn[62]), .inData_1(wireIn[63]), .outData_0(wireOut[62]), .outData_1(wireOut[63]), .ctrl(ctrl[31]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_32(.inData_0(wireIn[64]), .inData_1(wireIn[65]), .outData_0(wireOut[64]), .outData_1(wireOut[65]), .ctrl(ctrl[32]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_33(.inData_0(wireIn[66]), .inData_1(wireIn[67]), .outData_0(wireOut[66]), .outData_1(wireOut[67]), .ctrl(ctrl[33]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_34(.inData_0(wireIn[68]), .inData_1(wireIn[69]), .outData_0(wireOut[68]), .outData_1(wireOut[69]), .ctrl(ctrl[34]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_35(.inData_0(wireIn[70]), .inData_1(wireIn[71]), .outData_0(wireOut[70]), .outData_1(wireOut[71]), .ctrl(ctrl[35]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_36(.inData_0(wireIn[72]), .inData_1(wireIn[73]), .outData_0(wireOut[72]), .outData_1(wireOut[73]), .ctrl(ctrl[36]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_37(.inData_0(wireIn[74]), .inData_1(wireIn[75]), .outData_0(wireOut[74]), .outData_1(wireOut[75]), .ctrl(ctrl[37]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_38(.inData_0(wireIn[76]), .inData_1(wireIn[77]), .outData_0(wireOut[76]), .outData_1(wireOut[77]), .ctrl(ctrl[38]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_39(.inData_0(wireIn[78]), .inData_1(wireIn[79]), .outData_0(wireOut[78]), .outData_1(wireOut[79]), .ctrl(ctrl[39]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_40(.inData_0(wireIn[80]), .inData_1(wireIn[81]), .outData_0(wireOut[80]), .outData_1(wireOut[81]), .ctrl(ctrl[40]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_41(.inData_0(wireIn[82]), .inData_1(wireIn[83]), .outData_0(wireOut[82]), .outData_1(wireOut[83]), .ctrl(ctrl[41]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_42(.inData_0(wireIn[84]), .inData_1(wireIn[85]), .outData_0(wireOut[84]), .outData_1(wireOut[85]), .ctrl(ctrl[42]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_43(.inData_0(wireIn[86]), .inData_1(wireIn[87]), .outData_0(wireOut[86]), .outData_1(wireOut[87]), .ctrl(ctrl[43]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_44(.inData_0(wireIn[88]), .inData_1(wireIn[89]), .outData_0(wireOut[88]), .outData_1(wireOut[89]), .ctrl(ctrl[44]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_45(.inData_0(wireIn[90]), .inData_1(wireIn[91]), .outData_0(wireOut[90]), .outData_1(wireOut[91]), .ctrl(ctrl[45]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_46(.inData_0(wireIn[92]), .inData_1(wireIn[93]), .outData_0(wireOut[92]), .outData_1(wireOut[93]), .ctrl(ctrl[46]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_47(.inData_0(wireIn[94]), .inData_1(wireIn[95]), .outData_0(wireOut[94]), .outData_1(wireOut[95]), .ctrl(ctrl[47]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_48(.inData_0(wireIn[96]), .inData_1(wireIn[97]), .outData_0(wireOut[96]), .outData_1(wireOut[97]), .ctrl(ctrl[48]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_49(.inData_0(wireIn[98]), .inData_1(wireIn[99]), .outData_0(wireOut[98]), .outData_1(wireOut[99]), .ctrl(ctrl[49]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_50(.inData_0(wireIn[100]), .inData_1(wireIn[101]), .outData_0(wireOut[100]), .outData_1(wireOut[101]), .ctrl(ctrl[50]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_51(.inData_0(wireIn[102]), .inData_1(wireIn[103]), .outData_0(wireOut[102]), .outData_1(wireOut[103]), .ctrl(ctrl[51]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_52(.inData_0(wireIn[104]), .inData_1(wireIn[105]), .outData_0(wireOut[104]), .outData_1(wireOut[105]), .ctrl(ctrl[52]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_53(.inData_0(wireIn[106]), .inData_1(wireIn[107]), .outData_0(wireOut[106]), .outData_1(wireOut[107]), .ctrl(ctrl[53]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_54(.inData_0(wireIn[108]), .inData_1(wireIn[109]), .outData_0(wireOut[108]), .outData_1(wireOut[109]), .ctrl(ctrl[54]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_55(.inData_0(wireIn[110]), .inData_1(wireIn[111]), .outData_0(wireOut[110]), .outData_1(wireOut[111]), .ctrl(ctrl[55]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_56(.inData_0(wireIn[112]), .inData_1(wireIn[113]), .outData_0(wireOut[112]), .outData_1(wireOut[113]), .ctrl(ctrl[56]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_57(.inData_0(wireIn[114]), .inData_1(wireIn[115]), .outData_0(wireOut[114]), .outData_1(wireOut[115]), .ctrl(ctrl[57]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_58(.inData_0(wireIn[116]), .inData_1(wireIn[117]), .outData_0(wireOut[116]), .outData_1(wireOut[117]), .ctrl(ctrl[58]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_59(.inData_0(wireIn[118]), .inData_1(wireIn[119]), .outData_0(wireOut[118]), .outData_1(wireOut[119]), .ctrl(ctrl[59]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_60(.inData_0(wireIn[120]), .inData_1(wireIn[121]), .outData_0(wireOut[120]), .outData_1(wireOut[121]), .ctrl(ctrl[60]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_61(.inData_0(wireIn[122]), .inData_1(wireIn[123]), .outData_0(wireOut[122]), .outData_1(wireOut[123]), .ctrl(ctrl[61]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_62(.inData_0(wireIn[124]), .inData_1(wireIn[125]), .outData_0(wireOut[124]), .outData_1(wireOut[125]), .ctrl(ctrl[62]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_63(.inData_0(wireIn[126]), .inData_1(wireIn[127]), .outData_0(wireOut[126]), .outData_1(wireOut[127]), .ctrl(ctrl[63]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_64(.inData_0(wireIn[128]), .inData_1(wireIn[129]), .outData_0(wireOut[128]), .outData_1(wireOut[129]), .ctrl(ctrl[64]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_65(.inData_0(wireIn[130]), .inData_1(wireIn[131]), .outData_0(wireOut[130]), .outData_1(wireOut[131]), .ctrl(ctrl[65]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_66(.inData_0(wireIn[132]), .inData_1(wireIn[133]), .outData_0(wireOut[132]), .outData_1(wireOut[133]), .ctrl(ctrl[66]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_67(.inData_0(wireIn[134]), .inData_1(wireIn[135]), .outData_0(wireOut[134]), .outData_1(wireOut[135]), .ctrl(ctrl[67]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_68(.inData_0(wireIn[136]), .inData_1(wireIn[137]), .outData_0(wireOut[136]), .outData_1(wireOut[137]), .ctrl(ctrl[68]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_69(.inData_0(wireIn[138]), .inData_1(wireIn[139]), .outData_0(wireOut[138]), .outData_1(wireOut[139]), .ctrl(ctrl[69]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_70(.inData_0(wireIn[140]), .inData_1(wireIn[141]), .outData_0(wireOut[140]), .outData_1(wireOut[141]), .ctrl(ctrl[70]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_71(.inData_0(wireIn[142]), .inData_1(wireIn[143]), .outData_0(wireOut[142]), .outData_1(wireOut[143]), .ctrl(ctrl[71]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_72(.inData_0(wireIn[144]), .inData_1(wireIn[145]), .outData_0(wireOut[144]), .outData_1(wireOut[145]), .ctrl(ctrl[72]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_73(.inData_0(wireIn[146]), .inData_1(wireIn[147]), .outData_0(wireOut[146]), .outData_1(wireOut[147]), .ctrl(ctrl[73]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_74(.inData_0(wireIn[148]), .inData_1(wireIn[149]), .outData_0(wireOut[148]), .outData_1(wireOut[149]), .ctrl(ctrl[74]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_75(.inData_0(wireIn[150]), .inData_1(wireIn[151]), .outData_0(wireOut[150]), .outData_1(wireOut[151]), .ctrl(ctrl[75]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_76(.inData_0(wireIn[152]), .inData_1(wireIn[153]), .outData_0(wireOut[152]), .outData_1(wireOut[153]), .ctrl(ctrl[76]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_77(.inData_0(wireIn[154]), .inData_1(wireIn[155]), .outData_0(wireOut[154]), .outData_1(wireOut[155]), .ctrl(ctrl[77]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_78(.inData_0(wireIn[156]), .inData_1(wireIn[157]), .outData_0(wireOut[156]), .outData_1(wireOut[157]), .ctrl(ctrl[78]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_79(.inData_0(wireIn[158]), .inData_1(wireIn[159]), .outData_0(wireOut[158]), .outData_1(wireOut[159]), .ctrl(ctrl[79]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_80(.inData_0(wireIn[160]), .inData_1(wireIn[161]), .outData_0(wireOut[160]), .outData_1(wireOut[161]), .ctrl(ctrl[80]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_81(.inData_0(wireIn[162]), .inData_1(wireIn[163]), .outData_0(wireOut[162]), .outData_1(wireOut[163]), .ctrl(ctrl[81]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_82(.inData_0(wireIn[164]), .inData_1(wireIn[165]), .outData_0(wireOut[164]), .outData_1(wireOut[165]), .ctrl(ctrl[82]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_83(.inData_0(wireIn[166]), .inData_1(wireIn[167]), .outData_0(wireOut[166]), .outData_1(wireOut[167]), .ctrl(ctrl[83]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_84(.inData_0(wireIn[168]), .inData_1(wireIn[169]), .outData_0(wireOut[168]), .outData_1(wireOut[169]), .ctrl(ctrl[84]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_85(.inData_0(wireIn[170]), .inData_1(wireIn[171]), .outData_0(wireOut[170]), .outData_1(wireOut[171]), .ctrl(ctrl[85]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_86(.inData_0(wireIn[172]), .inData_1(wireIn[173]), .outData_0(wireOut[172]), .outData_1(wireOut[173]), .ctrl(ctrl[86]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_87(.inData_0(wireIn[174]), .inData_1(wireIn[175]), .outData_0(wireOut[174]), .outData_1(wireOut[175]), .ctrl(ctrl[87]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_88(.inData_0(wireIn[176]), .inData_1(wireIn[177]), .outData_0(wireOut[176]), .outData_1(wireOut[177]), .ctrl(ctrl[88]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_89(.inData_0(wireIn[178]), .inData_1(wireIn[179]), .outData_0(wireOut[178]), .outData_1(wireOut[179]), .ctrl(ctrl[89]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_90(.inData_0(wireIn[180]), .inData_1(wireIn[181]), .outData_0(wireOut[180]), .outData_1(wireOut[181]), .ctrl(ctrl[90]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_91(.inData_0(wireIn[182]), .inData_1(wireIn[183]), .outData_0(wireOut[182]), .outData_1(wireOut[183]), .ctrl(ctrl[91]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_92(.inData_0(wireIn[184]), .inData_1(wireIn[185]), .outData_0(wireOut[184]), .outData_1(wireOut[185]), .ctrl(ctrl[92]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_93(.inData_0(wireIn[186]), .inData_1(wireIn[187]), .outData_0(wireOut[186]), .outData_1(wireOut[187]), .ctrl(ctrl[93]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_94(.inData_0(wireIn[188]), .inData_1(wireIn[189]), .outData_0(wireOut[188]), .outData_1(wireOut[189]), .ctrl(ctrl[94]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_95(.inData_0(wireIn[190]), .inData_1(wireIn[191]), .outData_0(wireOut[190]), .outData_1(wireOut[191]), .ctrl(ctrl[95]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_96(.inData_0(wireIn[192]), .inData_1(wireIn[193]), .outData_0(wireOut[192]), .outData_1(wireOut[193]), .ctrl(ctrl[96]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_97(.inData_0(wireIn[194]), .inData_1(wireIn[195]), .outData_0(wireOut[194]), .outData_1(wireOut[195]), .ctrl(ctrl[97]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_98(.inData_0(wireIn[196]), .inData_1(wireIn[197]), .outData_0(wireOut[196]), .outData_1(wireOut[197]), .ctrl(ctrl[98]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_99(.inData_0(wireIn[198]), .inData_1(wireIn[199]), .outData_0(wireOut[198]), .outData_1(wireOut[199]), .ctrl(ctrl[99]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_100(.inData_0(wireIn[200]), .inData_1(wireIn[201]), .outData_0(wireOut[200]), .outData_1(wireOut[201]), .ctrl(ctrl[100]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_101(.inData_0(wireIn[202]), .inData_1(wireIn[203]), .outData_0(wireOut[202]), .outData_1(wireOut[203]), .ctrl(ctrl[101]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_102(.inData_0(wireIn[204]), .inData_1(wireIn[205]), .outData_0(wireOut[204]), .outData_1(wireOut[205]), .ctrl(ctrl[102]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_103(.inData_0(wireIn[206]), .inData_1(wireIn[207]), .outData_0(wireOut[206]), .outData_1(wireOut[207]), .ctrl(ctrl[103]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_104(.inData_0(wireIn[208]), .inData_1(wireIn[209]), .outData_0(wireOut[208]), .outData_1(wireOut[209]), .ctrl(ctrl[104]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_105(.inData_0(wireIn[210]), .inData_1(wireIn[211]), .outData_0(wireOut[210]), .outData_1(wireOut[211]), .ctrl(ctrl[105]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_106(.inData_0(wireIn[212]), .inData_1(wireIn[213]), .outData_0(wireOut[212]), .outData_1(wireOut[213]), .ctrl(ctrl[106]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_107(.inData_0(wireIn[214]), .inData_1(wireIn[215]), .outData_0(wireOut[214]), .outData_1(wireOut[215]), .ctrl(ctrl[107]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_108(.inData_0(wireIn[216]), .inData_1(wireIn[217]), .outData_0(wireOut[216]), .outData_1(wireOut[217]), .ctrl(ctrl[108]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_109(.inData_0(wireIn[218]), .inData_1(wireIn[219]), .outData_0(wireOut[218]), .outData_1(wireOut[219]), .ctrl(ctrl[109]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_110(.inData_0(wireIn[220]), .inData_1(wireIn[221]), .outData_0(wireOut[220]), .outData_1(wireOut[221]), .ctrl(ctrl[110]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_111(.inData_0(wireIn[222]), .inData_1(wireIn[223]), .outData_0(wireOut[222]), .outData_1(wireOut[223]), .ctrl(ctrl[111]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_112(.inData_0(wireIn[224]), .inData_1(wireIn[225]), .outData_0(wireOut[224]), .outData_1(wireOut[225]), .ctrl(ctrl[112]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_113(.inData_0(wireIn[226]), .inData_1(wireIn[227]), .outData_0(wireOut[226]), .outData_1(wireOut[227]), .ctrl(ctrl[113]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_114(.inData_0(wireIn[228]), .inData_1(wireIn[229]), .outData_0(wireOut[228]), .outData_1(wireOut[229]), .ctrl(ctrl[114]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_115(.inData_0(wireIn[230]), .inData_1(wireIn[231]), .outData_0(wireOut[230]), .outData_1(wireOut[231]), .ctrl(ctrl[115]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_116(.inData_0(wireIn[232]), .inData_1(wireIn[233]), .outData_0(wireOut[232]), .outData_1(wireOut[233]), .ctrl(ctrl[116]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_117(.inData_0(wireIn[234]), .inData_1(wireIn[235]), .outData_0(wireOut[234]), .outData_1(wireOut[235]), .ctrl(ctrl[117]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_118(.inData_0(wireIn[236]), .inData_1(wireIn[237]), .outData_0(wireOut[236]), .outData_1(wireOut[237]), .ctrl(ctrl[118]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_119(.inData_0(wireIn[238]), .inData_1(wireIn[239]), .outData_0(wireOut[238]), .outData_1(wireOut[239]), .ctrl(ctrl[119]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_120(.inData_0(wireIn[240]), .inData_1(wireIn[241]), .outData_0(wireOut[240]), .outData_1(wireOut[241]), .ctrl(ctrl[120]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_121(.inData_0(wireIn[242]), .inData_1(wireIn[243]), .outData_0(wireOut[242]), .outData_1(wireOut[243]), .ctrl(ctrl[121]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_122(.inData_0(wireIn[244]), .inData_1(wireIn[245]), .outData_0(wireOut[244]), .outData_1(wireOut[245]), .ctrl(ctrl[122]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_123(.inData_0(wireIn[246]), .inData_1(wireIn[247]), .outData_0(wireOut[246]), .outData_1(wireOut[247]), .ctrl(ctrl[123]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_124(.inData_0(wireIn[248]), .inData_1(wireIn[249]), .outData_0(wireOut[248]), .outData_1(wireOut[249]), .ctrl(ctrl[124]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_125(.inData_0(wireIn[250]), .inData_1(wireIn[251]), .outData_0(wireOut[250]), .outData_1(wireOut[251]), .ctrl(ctrl[125]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_126(.inData_0(wireIn[252]), .inData_1(wireIn[253]), .outData_0(wireOut[252]), .outData_1(wireOut[253]), .ctrl(ctrl[126]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_127(.inData_0(wireIn[254]), .inData_1(wireIn[255]), .outData_0(wireOut[254]), .outData_1(wireOut[255]), .ctrl(ctrl[127]), .clk(clk), .rst(rst));
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module wireCon_dp256_st5_L(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  assign wireOut[0] = wireIn[0];    
  assign wireOut[1] = wireIn[2];    
  assign wireOut[2] = wireIn[4];    
  assign wireOut[3] = wireIn[6];    
  assign wireOut[4] = wireIn[1];    
  assign wireOut[5] = wireIn[3];    
  assign wireOut[6] = wireIn[5];    
  assign wireOut[7] = wireIn[7];    
  assign wireOut[8] = wireIn[8];    
  assign wireOut[9] = wireIn[10];    
  assign wireOut[10] = wireIn[12];    
  assign wireOut[11] = wireIn[14];    
  assign wireOut[12] = wireIn[9];    
  assign wireOut[13] = wireIn[11];    
  assign wireOut[14] = wireIn[13];    
  assign wireOut[15] = wireIn[15];    
  assign wireOut[16] = wireIn[16];    
  assign wireOut[17] = wireIn[18];    
  assign wireOut[18] = wireIn[20];    
  assign wireOut[19] = wireIn[22];    
  assign wireOut[20] = wireIn[17];    
  assign wireOut[21] = wireIn[19];    
  assign wireOut[22] = wireIn[21];    
  assign wireOut[23] = wireIn[23];    
  assign wireOut[24] = wireIn[24];    
  assign wireOut[25] = wireIn[26];    
  assign wireOut[26] = wireIn[28];    
  assign wireOut[27] = wireIn[30];    
  assign wireOut[28] = wireIn[25];    
  assign wireOut[29] = wireIn[27];    
  assign wireOut[30] = wireIn[29];    
  assign wireOut[31] = wireIn[31];    
  assign wireOut[32] = wireIn[32];    
  assign wireOut[33] = wireIn[34];    
  assign wireOut[34] = wireIn[36];    
  assign wireOut[35] = wireIn[38];    
  assign wireOut[36] = wireIn[33];    
  assign wireOut[37] = wireIn[35];    
  assign wireOut[38] = wireIn[37];    
  assign wireOut[39] = wireIn[39];    
  assign wireOut[40] = wireIn[40];    
  assign wireOut[41] = wireIn[42];    
  assign wireOut[42] = wireIn[44];    
  assign wireOut[43] = wireIn[46];    
  assign wireOut[44] = wireIn[41];    
  assign wireOut[45] = wireIn[43];    
  assign wireOut[46] = wireIn[45];    
  assign wireOut[47] = wireIn[47];    
  assign wireOut[48] = wireIn[48];    
  assign wireOut[49] = wireIn[50];    
  assign wireOut[50] = wireIn[52];    
  assign wireOut[51] = wireIn[54];    
  assign wireOut[52] = wireIn[49];    
  assign wireOut[53] = wireIn[51];    
  assign wireOut[54] = wireIn[53];    
  assign wireOut[55] = wireIn[55];    
  assign wireOut[56] = wireIn[56];    
  assign wireOut[57] = wireIn[58];    
  assign wireOut[58] = wireIn[60];    
  assign wireOut[59] = wireIn[62];    
  assign wireOut[60] = wireIn[57];    
  assign wireOut[61] = wireIn[59];    
  assign wireOut[62] = wireIn[61];    
  assign wireOut[63] = wireIn[63];    
  assign wireOut[64] = wireIn[64];    
  assign wireOut[65] = wireIn[66];    
  assign wireOut[66] = wireIn[68];    
  assign wireOut[67] = wireIn[70];    
  assign wireOut[68] = wireIn[65];    
  assign wireOut[69] = wireIn[67];    
  assign wireOut[70] = wireIn[69];    
  assign wireOut[71] = wireIn[71];    
  assign wireOut[72] = wireIn[72];    
  assign wireOut[73] = wireIn[74];    
  assign wireOut[74] = wireIn[76];    
  assign wireOut[75] = wireIn[78];    
  assign wireOut[76] = wireIn[73];    
  assign wireOut[77] = wireIn[75];    
  assign wireOut[78] = wireIn[77];    
  assign wireOut[79] = wireIn[79];    
  assign wireOut[80] = wireIn[80];    
  assign wireOut[81] = wireIn[82];    
  assign wireOut[82] = wireIn[84];    
  assign wireOut[83] = wireIn[86];    
  assign wireOut[84] = wireIn[81];    
  assign wireOut[85] = wireIn[83];    
  assign wireOut[86] = wireIn[85];    
  assign wireOut[87] = wireIn[87];    
  assign wireOut[88] = wireIn[88];    
  assign wireOut[89] = wireIn[90];    
  assign wireOut[90] = wireIn[92];    
  assign wireOut[91] = wireIn[94];    
  assign wireOut[92] = wireIn[89];    
  assign wireOut[93] = wireIn[91];    
  assign wireOut[94] = wireIn[93];    
  assign wireOut[95] = wireIn[95];    
  assign wireOut[96] = wireIn[96];    
  assign wireOut[97] = wireIn[98];    
  assign wireOut[98] = wireIn[100];    
  assign wireOut[99] = wireIn[102];    
  assign wireOut[100] = wireIn[97];    
  assign wireOut[101] = wireIn[99];    
  assign wireOut[102] = wireIn[101];    
  assign wireOut[103] = wireIn[103];    
  assign wireOut[104] = wireIn[104];    
  assign wireOut[105] = wireIn[106];    
  assign wireOut[106] = wireIn[108];    
  assign wireOut[107] = wireIn[110];    
  assign wireOut[108] = wireIn[105];    
  assign wireOut[109] = wireIn[107];    
  assign wireOut[110] = wireIn[109];    
  assign wireOut[111] = wireIn[111];    
  assign wireOut[112] = wireIn[112];    
  assign wireOut[113] = wireIn[114];    
  assign wireOut[114] = wireIn[116];    
  assign wireOut[115] = wireIn[118];    
  assign wireOut[116] = wireIn[113];    
  assign wireOut[117] = wireIn[115];    
  assign wireOut[118] = wireIn[117];    
  assign wireOut[119] = wireIn[119];    
  assign wireOut[120] = wireIn[120];    
  assign wireOut[121] = wireIn[122];    
  assign wireOut[122] = wireIn[124];    
  assign wireOut[123] = wireIn[126];    
  assign wireOut[124] = wireIn[121];    
  assign wireOut[125] = wireIn[123];    
  assign wireOut[126] = wireIn[125];    
  assign wireOut[127] = wireIn[127];    
  assign wireOut[128] = wireIn[128];    
  assign wireOut[129] = wireIn[130];    
  assign wireOut[130] = wireIn[132];    
  assign wireOut[131] = wireIn[134];    
  assign wireOut[132] = wireIn[129];    
  assign wireOut[133] = wireIn[131];    
  assign wireOut[134] = wireIn[133];    
  assign wireOut[135] = wireIn[135];    
  assign wireOut[136] = wireIn[136];    
  assign wireOut[137] = wireIn[138];    
  assign wireOut[138] = wireIn[140];    
  assign wireOut[139] = wireIn[142];    
  assign wireOut[140] = wireIn[137];    
  assign wireOut[141] = wireIn[139];    
  assign wireOut[142] = wireIn[141];    
  assign wireOut[143] = wireIn[143];    
  assign wireOut[144] = wireIn[144];    
  assign wireOut[145] = wireIn[146];    
  assign wireOut[146] = wireIn[148];    
  assign wireOut[147] = wireIn[150];    
  assign wireOut[148] = wireIn[145];    
  assign wireOut[149] = wireIn[147];    
  assign wireOut[150] = wireIn[149];    
  assign wireOut[151] = wireIn[151];    
  assign wireOut[152] = wireIn[152];    
  assign wireOut[153] = wireIn[154];    
  assign wireOut[154] = wireIn[156];    
  assign wireOut[155] = wireIn[158];    
  assign wireOut[156] = wireIn[153];    
  assign wireOut[157] = wireIn[155];    
  assign wireOut[158] = wireIn[157];    
  assign wireOut[159] = wireIn[159];    
  assign wireOut[160] = wireIn[160];    
  assign wireOut[161] = wireIn[162];    
  assign wireOut[162] = wireIn[164];    
  assign wireOut[163] = wireIn[166];    
  assign wireOut[164] = wireIn[161];    
  assign wireOut[165] = wireIn[163];    
  assign wireOut[166] = wireIn[165];    
  assign wireOut[167] = wireIn[167];    
  assign wireOut[168] = wireIn[168];    
  assign wireOut[169] = wireIn[170];    
  assign wireOut[170] = wireIn[172];    
  assign wireOut[171] = wireIn[174];    
  assign wireOut[172] = wireIn[169];    
  assign wireOut[173] = wireIn[171];    
  assign wireOut[174] = wireIn[173];    
  assign wireOut[175] = wireIn[175];    
  assign wireOut[176] = wireIn[176];    
  assign wireOut[177] = wireIn[178];    
  assign wireOut[178] = wireIn[180];    
  assign wireOut[179] = wireIn[182];    
  assign wireOut[180] = wireIn[177];    
  assign wireOut[181] = wireIn[179];    
  assign wireOut[182] = wireIn[181];    
  assign wireOut[183] = wireIn[183];    
  assign wireOut[184] = wireIn[184];    
  assign wireOut[185] = wireIn[186];    
  assign wireOut[186] = wireIn[188];    
  assign wireOut[187] = wireIn[190];    
  assign wireOut[188] = wireIn[185];    
  assign wireOut[189] = wireIn[187];    
  assign wireOut[190] = wireIn[189];    
  assign wireOut[191] = wireIn[191];    
  assign wireOut[192] = wireIn[192];    
  assign wireOut[193] = wireIn[194];    
  assign wireOut[194] = wireIn[196];    
  assign wireOut[195] = wireIn[198];    
  assign wireOut[196] = wireIn[193];    
  assign wireOut[197] = wireIn[195];    
  assign wireOut[198] = wireIn[197];    
  assign wireOut[199] = wireIn[199];    
  assign wireOut[200] = wireIn[200];    
  assign wireOut[201] = wireIn[202];    
  assign wireOut[202] = wireIn[204];    
  assign wireOut[203] = wireIn[206];    
  assign wireOut[204] = wireIn[201];    
  assign wireOut[205] = wireIn[203];    
  assign wireOut[206] = wireIn[205];    
  assign wireOut[207] = wireIn[207];    
  assign wireOut[208] = wireIn[208];    
  assign wireOut[209] = wireIn[210];    
  assign wireOut[210] = wireIn[212];    
  assign wireOut[211] = wireIn[214];    
  assign wireOut[212] = wireIn[209];    
  assign wireOut[213] = wireIn[211];    
  assign wireOut[214] = wireIn[213];    
  assign wireOut[215] = wireIn[215];    
  assign wireOut[216] = wireIn[216];    
  assign wireOut[217] = wireIn[218];    
  assign wireOut[218] = wireIn[220];    
  assign wireOut[219] = wireIn[222];    
  assign wireOut[220] = wireIn[217];    
  assign wireOut[221] = wireIn[219];    
  assign wireOut[222] = wireIn[221];    
  assign wireOut[223] = wireIn[223];    
  assign wireOut[224] = wireIn[224];    
  assign wireOut[225] = wireIn[226];    
  assign wireOut[226] = wireIn[228];    
  assign wireOut[227] = wireIn[230];    
  assign wireOut[228] = wireIn[225];    
  assign wireOut[229] = wireIn[227];    
  assign wireOut[230] = wireIn[229];    
  assign wireOut[231] = wireIn[231];    
  assign wireOut[232] = wireIn[232];    
  assign wireOut[233] = wireIn[234];    
  assign wireOut[234] = wireIn[236];    
  assign wireOut[235] = wireIn[238];    
  assign wireOut[236] = wireIn[233];    
  assign wireOut[237] = wireIn[235];    
  assign wireOut[238] = wireIn[237];    
  assign wireOut[239] = wireIn[239];    
  assign wireOut[240] = wireIn[240];    
  assign wireOut[241] = wireIn[242];    
  assign wireOut[242] = wireIn[244];    
  assign wireOut[243] = wireIn[246];    
  assign wireOut[244] = wireIn[241];    
  assign wireOut[245] = wireIn[243];    
  assign wireOut[246] = wireIn[245];    
  assign wireOut[247] = wireIn[247];    
  assign wireOut[248] = wireIn[248];    
  assign wireOut[249] = wireIn[250];    
  assign wireOut[250] = wireIn[252];    
  assign wireOut[251] = wireIn[254];    
  assign wireOut[252] = wireIn[249];    
  assign wireOut[253] = wireIn[251];    
  assign wireOut[254] = wireIn[253];    
  assign wireOut[255] = wireIn[255];    
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module switches_stage_st6_0_L(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
ctrl,                            
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;                   
  input [128-1:0] ctrl;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  switch_2_2 switch_inst_0(.inData_0(wireIn[0]), .inData_1(wireIn[1]), .outData_0(wireOut[0]), .outData_1(wireOut[1]), .ctrl(ctrl[0]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_1(.inData_0(wireIn[2]), .inData_1(wireIn[3]), .outData_0(wireOut[2]), .outData_1(wireOut[3]), .ctrl(ctrl[1]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_2(.inData_0(wireIn[4]), .inData_1(wireIn[5]), .outData_0(wireOut[4]), .outData_1(wireOut[5]), .ctrl(ctrl[2]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_3(.inData_0(wireIn[6]), .inData_1(wireIn[7]), .outData_0(wireOut[6]), .outData_1(wireOut[7]), .ctrl(ctrl[3]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_4(.inData_0(wireIn[8]), .inData_1(wireIn[9]), .outData_0(wireOut[8]), .outData_1(wireOut[9]), .ctrl(ctrl[4]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_5(.inData_0(wireIn[10]), .inData_1(wireIn[11]), .outData_0(wireOut[10]), .outData_1(wireOut[11]), .ctrl(ctrl[5]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_6(.inData_0(wireIn[12]), .inData_1(wireIn[13]), .outData_0(wireOut[12]), .outData_1(wireOut[13]), .ctrl(ctrl[6]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_7(.inData_0(wireIn[14]), .inData_1(wireIn[15]), .outData_0(wireOut[14]), .outData_1(wireOut[15]), .ctrl(ctrl[7]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_8(.inData_0(wireIn[16]), .inData_1(wireIn[17]), .outData_0(wireOut[16]), .outData_1(wireOut[17]), .ctrl(ctrl[8]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_9(.inData_0(wireIn[18]), .inData_1(wireIn[19]), .outData_0(wireOut[18]), .outData_1(wireOut[19]), .ctrl(ctrl[9]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_10(.inData_0(wireIn[20]), .inData_1(wireIn[21]), .outData_0(wireOut[20]), .outData_1(wireOut[21]), .ctrl(ctrl[10]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_11(.inData_0(wireIn[22]), .inData_1(wireIn[23]), .outData_0(wireOut[22]), .outData_1(wireOut[23]), .ctrl(ctrl[11]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_12(.inData_0(wireIn[24]), .inData_1(wireIn[25]), .outData_0(wireOut[24]), .outData_1(wireOut[25]), .ctrl(ctrl[12]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_13(.inData_0(wireIn[26]), .inData_1(wireIn[27]), .outData_0(wireOut[26]), .outData_1(wireOut[27]), .ctrl(ctrl[13]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_14(.inData_0(wireIn[28]), .inData_1(wireIn[29]), .outData_0(wireOut[28]), .outData_1(wireOut[29]), .ctrl(ctrl[14]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_15(.inData_0(wireIn[30]), .inData_1(wireIn[31]), .outData_0(wireOut[30]), .outData_1(wireOut[31]), .ctrl(ctrl[15]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_16(.inData_0(wireIn[32]), .inData_1(wireIn[33]), .outData_0(wireOut[32]), .outData_1(wireOut[33]), .ctrl(ctrl[16]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_17(.inData_0(wireIn[34]), .inData_1(wireIn[35]), .outData_0(wireOut[34]), .outData_1(wireOut[35]), .ctrl(ctrl[17]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_18(.inData_0(wireIn[36]), .inData_1(wireIn[37]), .outData_0(wireOut[36]), .outData_1(wireOut[37]), .ctrl(ctrl[18]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_19(.inData_0(wireIn[38]), .inData_1(wireIn[39]), .outData_0(wireOut[38]), .outData_1(wireOut[39]), .ctrl(ctrl[19]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_20(.inData_0(wireIn[40]), .inData_1(wireIn[41]), .outData_0(wireOut[40]), .outData_1(wireOut[41]), .ctrl(ctrl[20]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_21(.inData_0(wireIn[42]), .inData_1(wireIn[43]), .outData_0(wireOut[42]), .outData_1(wireOut[43]), .ctrl(ctrl[21]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_22(.inData_0(wireIn[44]), .inData_1(wireIn[45]), .outData_0(wireOut[44]), .outData_1(wireOut[45]), .ctrl(ctrl[22]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_23(.inData_0(wireIn[46]), .inData_1(wireIn[47]), .outData_0(wireOut[46]), .outData_1(wireOut[47]), .ctrl(ctrl[23]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_24(.inData_0(wireIn[48]), .inData_1(wireIn[49]), .outData_0(wireOut[48]), .outData_1(wireOut[49]), .ctrl(ctrl[24]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_25(.inData_0(wireIn[50]), .inData_1(wireIn[51]), .outData_0(wireOut[50]), .outData_1(wireOut[51]), .ctrl(ctrl[25]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_26(.inData_0(wireIn[52]), .inData_1(wireIn[53]), .outData_0(wireOut[52]), .outData_1(wireOut[53]), .ctrl(ctrl[26]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_27(.inData_0(wireIn[54]), .inData_1(wireIn[55]), .outData_0(wireOut[54]), .outData_1(wireOut[55]), .ctrl(ctrl[27]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_28(.inData_0(wireIn[56]), .inData_1(wireIn[57]), .outData_0(wireOut[56]), .outData_1(wireOut[57]), .ctrl(ctrl[28]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_29(.inData_0(wireIn[58]), .inData_1(wireIn[59]), .outData_0(wireOut[58]), .outData_1(wireOut[59]), .ctrl(ctrl[29]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_30(.inData_0(wireIn[60]), .inData_1(wireIn[61]), .outData_0(wireOut[60]), .outData_1(wireOut[61]), .ctrl(ctrl[30]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_31(.inData_0(wireIn[62]), .inData_1(wireIn[63]), .outData_0(wireOut[62]), .outData_1(wireOut[63]), .ctrl(ctrl[31]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_32(.inData_0(wireIn[64]), .inData_1(wireIn[65]), .outData_0(wireOut[64]), .outData_1(wireOut[65]), .ctrl(ctrl[32]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_33(.inData_0(wireIn[66]), .inData_1(wireIn[67]), .outData_0(wireOut[66]), .outData_1(wireOut[67]), .ctrl(ctrl[33]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_34(.inData_0(wireIn[68]), .inData_1(wireIn[69]), .outData_0(wireOut[68]), .outData_1(wireOut[69]), .ctrl(ctrl[34]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_35(.inData_0(wireIn[70]), .inData_1(wireIn[71]), .outData_0(wireOut[70]), .outData_1(wireOut[71]), .ctrl(ctrl[35]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_36(.inData_0(wireIn[72]), .inData_1(wireIn[73]), .outData_0(wireOut[72]), .outData_1(wireOut[73]), .ctrl(ctrl[36]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_37(.inData_0(wireIn[74]), .inData_1(wireIn[75]), .outData_0(wireOut[74]), .outData_1(wireOut[75]), .ctrl(ctrl[37]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_38(.inData_0(wireIn[76]), .inData_1(wireIn[77]), .outData_0(wireOut[76]), .outData_1(wireOut[77]), .ctrl(ctrl[38]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_39(.inData_0(wireIn[78]), .inData_1(wireIn[79]), .outData_0(wireOut[78]), .outData_1(wireOut[79]), .ctrl(ctrl[39]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_40(.inData_0(wireIn[80]), .inData_1(wireIn[81]), .outData_0(wireOut[80]), .outData_1(wireOut[81]), .ctrl(ctrl[40]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_41(.inData_0(wireIn[82]), .inData_1(wireIn[83]), .outData_0(wireOut[82]), .outData_1(wireOut[83]), .ctrl(ctrl[41]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_42(.inData_0(wireIn[84]), .inData_1(wireIn[85]), .outData_0(wireOut[84]), .outData_1(wireOut[85]), .ctrl(ctrl[42]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_43(.inData_0(wireIn[86]), .inData_1(wireIn[87]), .outData_0(wireOut[86]), .outData_1(wireOut[87]), .ctrl(ctrl[43]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_44(.inData_0(wireIn[88]), .inData_1(wireIn[89]), .outData_0(wireOut[88]), .outData_1(wireOut[89]), .ctrl(ctrl[44]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_45(.inData_0(wireIn[90]), .inData_1(wireIn[91]), .outData_0(wireOut[90]), .outData_1(wireOut[91]), .ctrl(ctrl[45]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_46(.inData_0(wireIn[92]), .inData_1(wireIn[93]), .outData_0(wireOut[92]), .outData_1(wireOut[93]), .ctrl(ctrl[46]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_47(.inData_0(wireIn[94]), .inData_1(wireIn[95]), .outData_0(wireOut[94]), .outData_1(wireOut[95]), .ctrl(ctrl[47]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_48(.inData_0(wireIn[96]), .inData_1(wireIn[97]), .outData_0(wireOut[96]), .outData_1(wireOut[97]), .ctrl(ctrl[48]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_49(.inData_0(wireIn[98]), .inData_1(wireIn[99]), .outData_0(wireOut[98]), .outData_1(wireOut[99]), .ctrl(ctrl[49]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_50(.inData_0(wireIn[100]), .inData_1(wireIn[101]), .outData_0(wireOut[100]), .outData_1(wireOut[101]), .ctrl(ctrl[50]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_51(.inData_0(wireIn[102]), .inData_1(wireIn[103]), .outData_0(wireOut[102]), .outData_1(wireOut[103]), .ctrl(ctrl[51]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_52(.inData_0(wireIn[104]), .inData_1(wireIn[105]), .outData_0(wireOut[104]), .outData_1(wireOut[105]), .ctrl(ctrl[52]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_53(.inData_0(wireIn[106]), .inData_1(wireIn[107]), .outData_0(wireOut[106]), .outData_1(wireOut[107]), .ctrl(ctrl[53]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_54(.inData_0(wireIn[108]), .inData_1(wireIn[109]), .outData_0(wireOut[108]), .outData_1(wireOut[109]), .ctrl(ctrl[54]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_55(.inData_0(wireIn[110]), .inData_1(wireIn[111]), .outData_0(wireOut[110]), .outData_1(wireOut[111]), .ctrl(ctrl[55]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_56(.inData_0(wireIn[112]), .inData_1(wireIn[113]), .outData_0(wireOut[112]), .outData_1(wireOut[113]), .ctrl(ctrl[56]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_57(.inData_0(wireIn[114]), .inData_1(wireIn[115]), .outData_0(wireOut[114]), .outData_1(wireOut[115]), .ctrl(ctrl[57]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_58(.inData_0(wireIn[116]), .inData_1(wireIn[117]), .outData_0(wireOut[116]), .outData_1(wireOut[117]), .ctrl(ctrl[58]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_59(.inData_0(wireIn[118]), .inData_1(wireIn[119]), .outData_0(wireOut[118]), .outData_1(wireOut[119]), .ctrl(ctrl[59]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_60(.inData_0(wireIn[120]), .inData_1(wireIn[121]), .outData_0(wireOut[120]), .outData_1(wireOut[121]), .ctrl(ctrl[60]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_61(.inData_0(wireIn[122]), .inData_1(wireIn[123]), .outData_0(wireOut[122]), .outData_1(wireOut[123]), .ctrl(ctrl[61]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_62(.inData_0(wireIn[124]), .inData_1(wireIn[125]), .outData_0(wireOut[124]), .outData_1(wireOut[125]), .ctrl(ctrl[62]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_63(.inData_0(wireIn[126]), .inData_1(wireIn[127]), .outData_0(wireOut[126]), .outData_1(wireOut[127]), .ctrl(ctrl[63]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_64(.inData_0(wireIn[128]), .inData_1(wireIn[129]), .outData_0(wireOut[128]), .outData_1(wireOut[129]), .ctrl(ctrl[64]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_65(.inData_0(wireIn[130]), .inData_1(wireIn[131]), .outData_0(wireOut[130]), .outData_1(wireOut[131]), .ctrl(ctrl[65]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_66(.inData_0(wireIn[132]), .inData_1(wireIn[133]), .outData_0(wireOut[132]), .outData_1(wireOut[133]), .ctrl(ctrl[66]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_67(.inData_0(wireIn[134]), .inData_1(wireIn[135]), .outData_0(wireOut[134]), .outData_1(wireOut[135]), .ctrl(ctrl[67]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_68(.inData_0(wireIn[136]), .inData_1(wireIn[137]), .outData_0(wireOut[136]), .outData_1(wireOut[137]), .ctrl(ctrl[68]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_69(.inData_0(wireIn[138]), .inData_1(wireIn[139]), .outData_0(wireOut[138]), .outData_1(wireOut[139]), .ctrl(ctrl[69]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_70(.inData_0(wireIn[140]), .inData_1(wireIn[141]), .outData_0(wireOut[140]), .outData_1(wireOut[141]), .ctrl(ctrl[70]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_71(.inData_0(wireIn[142]), .inData_1(wireIn[143]), .outData_0(wireOut[142]), .outData_1(wireOut[143]), .ctrl(ctrl[71]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_72(.inData_0(wireIn[144]), .inData_1(wireIn[145]), .outData_0(wireOut[144]), .outData_1(wireOut[145]), .ctrl(ctrl[72]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_73(.inData_0(wireIn[146]), .inData_1(wireIn[147]), .outData_0(wireOut[146]), .outData_1(wireOut[147]), .ctrl(ctrl[73]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_74(.inData_0(wireIn[148]), .inData_1(wireIn[149]), .outData_0(wireOut[148]), .outData_1(wireOut[149]), .ctrl(ctrl[74]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_75(.inData_0(wireIn[150]), .inData_1(wireIn[151]), .outData_0(wireOut[150]), .outData_1(wireOut[151]), .ctrl(ctrl[75]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_76(.inData_0(wireIn[152]), .inData_1(wireIn[153]), .outData_0(wireOut[152]), .outData_1(wireOut[153]), .ctrl(ctrl[76]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_77(.inData_0(wireIn[154]), .inData_1(wireIn[155]), .outData_0(wireOut[154]), .outData_1(wireOut[155]), .ctrl(ctrl[77]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_78(.inData_0(wireIn[156]), .inData_1(wireIn[157]), .outData_0(wireOut[156]), .outData_1(wireOut[157]), .ctrl(ctrl[78]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_79(.inData_0(wireIn[158]), .inData_1(wireIn[159]), .outData_0(wireOut[158]), .outData_1(wireOut[159]), .ctrl(ctrl[79]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_80(.inData_0(wireIn[160]), .inData_1(wireIn[161]), .outData_0(wireOut[160]), .outData_1(wireOut[161]), .ctrl(ctrl[80]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_81(.inData_0(wireIn[162]), .inData_1(wireIn[163]), .outData_0(wireOut[162]), .outData_1(wireOut[163]), .ctrl(ctrl[81]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_82(.inData_0(wireIn[164]), .inData_1(wireIn[165]), .outData_0(wireOut[164]), .outData_1(wireOut[165]), .ctrl(ctrl[82]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_83(.inData_0(wireIn[166]), .inData_1(wireIn[167]), .outData_0(wireOut[166]), .outData_1(wireOut[167]), .ctrl(ctrl[83]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_84(.inData_0(wireIn[168]), .inData_1(wireIn[169]), .outData_0(wireOut[168]), .outData_1(wireOut[169]), .ctrl(ctrl[84]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_85(.inData_0(wireIn[170]), .inData_1(wireIn[171]), .outData_0(wireOut[170]), .outData_1(wireOut[171]), .ctrl(ctrl[85]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_86(.inData_0(wireIn[172]), .inData_1(wireIn[173]), .outData_0(wireOut[172]), .outData_1(wireOut[173]), .ctrl(ctrl[86]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_87(.inData_0(wireIn[174]), .inData_1(wireIn[175]), .outData_0(wireOut[174]), .outData_1(wireOut[175]), .ctrl(ctrl[87]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_88(.inData_0(wireIn[176]), .inData_1(wireIn[177]), .outData_0(wireOut[176]), .outData_1(wireOut[177]), .ctrl(ctrl[88]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_89(.inData_0(wireIn[178]), .inData_1(wireIn[179]), .outData_0(wireOut[178]), .outData_1(wireOut[179]), .ctrl(ctrl[89]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_90(.inData_0(wireIn[180]), .inData_1(wireIn[181]), .outData_0(wireOut[180]), .outData_1(wireOut[181]), .ctrl(ctrl[90]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_91(.inData_0(wireIn[182]), .inData_1(wireIn[183]), .outData_0(wireOut[182]), .outData_1(wireOut[183]), .ctrl(ctrl[91]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_92(.inData_0(wireIn[184]), .inData_1(wireIn[185]), .outData_0(wireOut[184]), .outData_1(wireOut[185]), .ctrl(ctrl[92]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_93(.inData_0(wireIn[186]), .inData_1(wireIn[187]), .outData_0(wireOut[186]), .outData_1(wireOut[187]), .ctrl(ctrl[93]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_94(.inData_0(wireIn[188]), .inData_1(wireIn[189]), .outData_0(wireOut[188]), .outData_1(wireOut[189]), .ctrl(ctrl[94]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_95(.inData_0(wireIn[190]), .inData_1(wireIn[191]), .outData_0(wireOut[190]), .outData_1(wireOut[191]), .ctrl(ctrl[95]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_96(.inData_0(wireIn[192]), .inData_1(wireIn[193]), .outData_0(wireOut[192]), .outData_1(wireOut[193]), .ctrl(ctrl[96]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_97(.inData_0(wireIn[194]), .inData_1(wireIn[195]), .outData_0(wireOut[194]), .outData_1(wireOut[195]), .ctrl(ctrl[97]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_98(.inData_0(wireIn[196]), .inData_1(wireIn[197]), .outData_0(wireOut[196]), .outData_1(wireOut[197]), .ctrl(ctrl[98]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_99(.inData_0(wireIn[198]), .inData_1(wireIn[199]), .outData_0(wireOut[198]), .outData_1(wireOut[199]), .ctrl(ctrl[99]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_100(.inData_0(wireIn[200]), .inData_1(wireIn[201]), .outData_0(wireOut[200]), .outData_1(wireOut[201]), .ctrl(ctrl[100]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_101(.inData_0(wireIn[202]), .inData_1(wireIn[203]), .outData_0(wireOut[202]), .outData_1(wireOut[203]), .ctrl(ctrl[101]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_102(.inData_0(wireIn[204]), .inData_1(wireIn[205]), .outData_0(wireOut[204]), .outData_1(wireOut[205]), .ctrl(ctrl[102]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_103(.inData_0(wireIn[206]), .inData_1(wireIn[207]), .outData_0(wireOut[206]), .outData_1(wireOut[207]), .ctrl(ctrl[103]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_104(.inData_0(wireIn[208]), .inData_1(wireIn[209]), .outData_0(wireOut[208]), .outData_1(wireOut[209]), .ctrl(ctrl[104]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_105(.inData_0(wireIn[210]), .inData_1(wireIn[211]), .outData_0(wireOut[210]), .outData_1(wireOut[211]), .ctrl(ctrl[105]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_106(.inData_0(wireIn[212]), .inData_1(wireIn[213]), .outData_0(wireOut[212]), .outData_1(wireOut[213]), .ctrl(ctrl[106]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_107(.inData_0(wireIn[214]), .inData_1(wireIn[215]), .outData_0(wireOut[214]), .outData_1(wireOut[215]), .ctrl(ctrl[107]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_108(.inData_0(wireIn[216]), .inData_1(wireIn[217]), .outData_0(wireOut[216]), .outData_1(wireOut[217]), .ctrl(ctrl[108]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_109(.inData_0(wireIn[218]), .inData_1(wireIn[219]), .outData_0(wireOut[218]), .outData_1(wireOut[219]), .ctrl(ctrl[109]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_110(.inData_0(wireIn[220]), .inData_1(wireIn[221]), .outData_0(wireOut[220]), .outData_1(wireOut[221]), .ctrl(ctrl[110]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_111(.inData_0(wireIn[222]), .inData_1(wireIn[223]), .outData_0(wireOut[222]), .outData_1(wireOut[223]), .ctrl(ctrl[111]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_112(.inData_0(wireIn[224]), .inData_1(wireIn[225]), .outData_0(wireOut[224]), .outData_1(wireOut[225]), .ctrl(ctrl[112]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_113(.inData_0(wireIn[226]), .inData_1(wireIn[227]), .outData_0(wireOut[226]), .outData_1(wireOut[227]), .ctrl(ctrl[113]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_114(.inData_0(wireIn[228]), .inData_1(wireIn[229]), .outData_0(wireOut[228]), .outData_1(wireOut[229]), .ctrl(ctrl[114]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_115(.inData_0(wireIn[230]), .inData_1(wireIn[231]), .outData_0(wireOut[230]), .outData_1(wireOut[231]), .ctrl(ctrl[115]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_116(.inData_0(wireIn[232]), .inData_1(wireIn[233]), .outData_0(wireOut[232]), .outData_1(wireOut[233]), .ctrl(ctrl[116]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_117(.inData_0(wireIn[234]), .inData_1(wireIn[235]), .outData_0(wireOut[234]), .outData_1(wireOut[235]), .ctrl(ctrl[117]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_118(.inData_0(wireIn[236]), .inData_1(wireIn[237]), .outData_0(wireOut[236]), .outData_1(wireOut[237]), .ctrl(ctrl[118]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_119(.inData_0(wireIn[238]), .inData_1(wireIn[239]), .outData_0(wireOut[238]), .outData_1(wireOut[239]), .ctrl(ctrl[119]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_120(.inData_0(wireIn[240]), .inData_1(wireIn[241]), .outData_0(wireOut[240]), .outData_1(wireOut[241]), .ctrl(ctrl[120]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_121(.inData_0(wireIn[242]), .inData_1(wireIn[243]), .outData_0(wireOut[242]), .outData_1(wireOut[243]), .ctrl(ctrl[121]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_122(.inData_0(wireIn[244]), .inData_1(wireIn[245]), .outData_0(wireOut[244]), .outData_1(wireOut[245]), .ctrl(ctrl[122]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_123(.inData_0(wireIn[246]), .inData_1(wireIn[247]), .outData_0(wireOut[246]), .outData_1(wireOut[247]), .ctrl(ctrl[123]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_124(.inData_0(wireIn[248]), .inData_1(wireIn[249]), .outData_0(wireOut[248]), .outData_1(wireOut[249]), .ctrl(ctrl[124]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_125(.inData_0(wireIn[250]), .inData_1(wireIn[251]), .outData_0(wireOut[250]), .outData_1(wireOut[251]), .ctrl(ctrl[125]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_126(.inData_0(wireIn[252]), .inData_1(wireIn[253]), .outData_0(wireOut[252]), .outData_1(wireOut[253]), .ctrl(ctrl[126]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_127(.inData_0(wireIn[254]), .inData_1(wireIn[255]), .outData_0(wireOut[254]), .outData_1(wireOut[255]), .ctrl(ctrl[127]), .clk(clk), .rst(rst));
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module wireCon_dp256_st6_L(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  assign wireOut[0] = wireIn[0];    
  assign wireOut[1] = wireIn[2];    
  assign wireOut[2] = wireIn[1];    
  assign wireOut[3] = wireIn[3];    
  assign wireOut[4] = wireIn[4];    
  assign wireOut[5] = wireIn[6];    
  assign wireOut[6] = wireIn[5];    
  assign wireOut[7] = wireIn[7];    
  assign wireOut[8] = wireIn[8];    
  assign wireOut[9] = wireIn[10];    
  assign wireOut[10] = wireIn[9];    
  assign wireOut[11] = wireIn[11];    
  assign wireOut[12] = wireIn[12];    
  assign wireOut[13] = wireIn[14];    
  assign wireOut[14] = wireIn[13];    
  assign wireOut[15] = wireIn[15];    
  assign wireOut[16] = wireIn[16];    
  assign wireOut[17] = wireIn[18];    
  assign wireOut[18] = wireIn[17];    
  assign wireOut[19] = wireIn[19];    
  assign wireOut[20] = wireIn[20];    
  assign wireOut[21] = wireIn[22];    
  assign wireOut[22] = wireIn[21];    
  assign wireOut[23] = wireIn[23];    
  assign wireOut[24] = wireIn[24];    
  assign wireOut[25] = wireIn[26];    
  assign wireOut[26] = wireIn[25];    
  assign wireOut[27] = wireIn[27];    
  assign wireOut[28] = wireIn[28];    
  assign wireOut[29] = wireIn[30];    
  assign wireOut[30] = wireIn[29];    
  assign wireOut[31] = wireIn[31];    
  assign wireOut[32] = wireIn[32];    
  assign wireOut[33] = wireIn[34];    
  assign wireOut[34] = wireIn[33];    
  assign wireOut[35] = wireIn[35];    
  assign wireOut[36] = wireIn[36];    
  assign wireOut[37] = wireIn[38];    
  assign wireOut[38] = wireIn[37];    
  assign wireOut[39] = wireIn[39];    
  assign wireOut[40] = wireIn[40];    
  assign wireOut[41] = wireIn[42];    
  assign wireOut[42] = wireIn[41];    
  assign wireOut[43] = wireIn[43];    
  assign wireOut[44] = wireIn[44];    
  assign wireOut[45] = wireIn[46];    
  assign wireOut[46] = wireIn[45];    
  assign wireOut[47] = wireIn[47];    
  assign wireOut[48] = wireIn[48];    
  assign wireOut[49] = wireIn[50];    
  assign wireOut[50] = wireIn[49];    
  assign wireOut[51] = wireIn[51];    
  assign wireOut[52] = wireIn[52];    
  assign wireOut[53] = wireIn[54];    
  assign wireOut[54] = wireIn[53];    
  assign wireOut[55] = wireIn[55];    
  assign wireOut[56] = wireIn[56];    
  assign wireOut[57] = wireIn[58];    
  assign wireOut[58] = wireIn[57];    
  assign wireOut[59] = wireIn[59];    
  assign wireOut[60] = wireIn[60];    
  assign wireOut[61] = wireIn[62];    
  assign wireOut[62] = wireIn[61];    
  assign wireOut[63] = wireIn[63];    
  assign wireOut[64] = wireIn[64];    
  assign wireOut[65] = wireIn[66];    
  assign wireOut[66] = wireIn[65];    
  assign wireOut[67] = wireIn[67];    
  assign wireOut[68] = wireIn[68];    
  assign wireOut[69] = wireIn[70];    
  assign wireOut[70] = wireIn[69];    
  assign wireOut[71] = wireIn[71];    
  assign wireOut[72] = wireIn[72];    
  assign wireOut[73] = wireIn[74];    
  assign wireOut[74] = wireIn[73];    
  assign wireOut[75] = wireIn[75];    
  assign wireOut[76] = wireIn[76];    
  assign wireOut[77] = wireIn[78];    
  assign wireOut[78] = wireIn[77];    
  assign wireOut[79] = wireIn[79];    
  assign wireOut[80] = wireIn[80];    
  assign wireOut[81] = wireIn[82];    
  assign wireOut[82] = wireIn[81];    
  assign wireOut[83] = wireIn[83];    
  assign wireOut[84] = wireIn[84];    
  assign wireOut[85] = wireIn[86];    
  assign wireOut[86] = wireIn[85];    
  assign wireOut[87] = wireIn[87];    
  assign wireOut[88] = wireIn[88];    
  assign wireOut[89] = wireIn[90];    
  assign wireOut[90] = wireIn[89];    
  assign wireOut[91] = wireIn[91];    
  assign wireOut[92] = wireIn[92];    
  assign wireOut[93] = wireIn[94];    
  assign wireOut[94] = wireIn[93];    
  assign wireOut[95] = wireIn[95];    
  assign wireOut[96] = wireIn[96];    
  assign wireOut[97] = wireIn[98];    
  assign wireOut[98] = wireIn[97];    
  assign wireOut[99] = wireIn[99];    
  assign wireOut[100] = wireIn[100];    
  assign wireOut[101] = wireIn[102];    
  assign wireOut[102] = wireIn[101];    
  assign wireOut[103] = wireIn[103];    
  assign wireOut[104] = wireIn[104];    
  assign wireOut[105] = wireIn[106];    
  assign wireOut[106] = wireIn[105];    
  assign wireOut[107] = wireIn[107];    
  assign wireOut[108] = wireIn[108];    
  assign wireOut[109] = wireIn[110];    
  assign wireOut[110] = wireIn[109];    
  assign wireOut[111] = wireIn[111];    
  assign wireOut[112] = wireIn[112];    
  assign wireOut[113] = wireIn[114];    
  assign wireOut[114] = wireIn[113];    
  assign wireOut[115] = wireIn[115];    
  assign wireOut[116] = wireIn[116];    
  assign wireOut[117] = wireIn[118];    
  assign wireOut[118] = wireIn[117];    
  assign wireOut[119] = wireIn[119];    
  assign wireOut[120] = wireIn[120];    
  assign wireOut[121] = wireIn[122];    
  assign wireOut[122] = wireIn[121];    
  assign wireOut[123] = wireIn[123];    
  assign wireOut[124] = wireIn[124];    
  assign wireOut[125] = wireIn[126];    
  assign wireOut[126] = wireIn[125];    
  assign wireOut[127] = wireIn[127];    
  assign wireOut[128] = wireIn[128];    
  assign wireOut[129] = wireIn[130];    
  assign wireOut[130] = wireIn[129];    
  assign wireOut[131] = wireIn[131];    
  assign wireOut[132] = wireIn[132];    
  assign wireOut[133] = wireIn[134];    
  assign wireOut[134] = wireIn[133];    
  assign wireOut[135] = wireIn[135];    
  assign wireOut[136] = wireIn[136];    
  assign wireOut[137] = wireIn[138];    
  assign wireOut[138] = wireIn[137];    
  assign wireOut[139] = wireIn[139];    
  assign wireOut[140] = wireIn[140];    
  assign wireOut[141] = wireIn[142];    
  assign wireOut[142] = wireIn[141];    
  assign wireOut[143] = wireIn[143];    
  assign wireOut[144] = wireIn[144];    
  assign wireOut[145] = wireIn[146];    
  assign wireOut[146] = wireIn[145];    
  assign wireOut[147] = wireIn[147];    
  assign wireOut[148] = wireIn[148];    
  assign wireOut[149] = wireIn[150];    
  assign wireOut[150] = wireIn[149];    
  assign wireOut[151] = wireIn[151];    
  assign wireOut[152] = wireIn[152];    
  assign wireOut[153] = wireIn[154];    
  assign wireOut[154] = wireIn[153];    
  assign wireOut[155] = wireIn[155];    
  assign wireOut[156] = wireIn[156];    
  assign wireOut[157] = wireIn[158];    
  assign wireOut[158] = wireIn[157];    
  assign wireOut[159] = wireIn[159];    
  assign wireOut[160] = wireIn[160];    
  assign wireOut[161] = wireIn[162];    
  assign wireOut[162] = wireIn[161];    
  assign wireOut[163] = wireIn[163];    
  assign wireOut[164] = wireIn[164];    
  assign wireOut[165] = wireIn[166];    
  assign wireOut[166] = wireIn[165];    
  assign wireOut[167] = wireIn[167];    
  assign wireOut[168] = wireIn[168];    
  assign wireOut[169] = wireIn[170];    
  assign wireOut[170] = wireIn[169];    
  assign wireOut[171] = wireIn[171];    
  assign wireOut[172] = wireIn[172];    
  assign wireOut[173] = wireIn[174];    
  assign wireOut[174] = wireIn[173];    
  assign wireOut[175] = wireIn[175];    
  assign wireOut[176] = wireIn[176];    
  assign wireOut[177] = wireIn[178];    
  assign wireOut[178] = wireIn[177];    
  assign wireOut[179] = wireIn[179];    
  assign wireOut[180] = wireIn[180];    
  assign wireOut[181] = wireIn[182];    
  assign wireOut[182] = wireIn[181];    
  assign wireOut[183] = wireIn[183];    
  assign wireOut[184] = wireIn[184];    
  assign wireOut[185] = wireIn[186];    
  assign wireOut[186] = wireIn[185];    
  assign wireOut[187] = wireIn[187];    
  assign wireOut[188] = wireIn[188];    
  assign wireOut[189] = wireIn[190];    
  assign wireOut[190] = wireIn[189];    
  assign wireOut[191] = wireIn[191];    
  assign wireOut[192] = wireIn[192];    
  assign wireOut[193] = wireIn[194];    
  assign wireOut[194] = wireIn[193];    
  assign wireOut[195] = wireIn[195];    
  assign wireOut[196] = wireIn[196];    
  assign wireOut[197] = wireIn[198];    
  assign wireOut[198] = wireIn[197];    
  assign wireOut[199] = wireIn[199];    
  assign wireOut[200] = wireIn[200];    
  assign wireOut[201] = wireIn[202];    
  assign wireOut[202] = wireIn[201];    
  assign wireOut[203] = wireIn[203];    
  assign wireOut[204] = wireIn[204];    
  assign wireOut[205] = wireIn[206];    
  assign wireOut[206] = wireIn[205];    
  assign wireOut[207] = wireIn[207];    
  assign wireOut[208] = wireIn[208];    
  assign wireOut[209] = wireIn[210];    
  assign wireOut[210] = wireIn[209];    
  assign wireOut[211] = wireIn[211];    
  assign wireOut[212] = wireIn[212];    
  assign wireOut[213] = wireIn[214];    
  assign wireOut[214] = wireIn[213];    
  assign wireOut[215] = wireIn[215];    
  assign wireOut[216] = wireIn[216];    
  assign wireOut[217] = wireIn[218];    
  assign wireOut[218] = wireIn[217];    
  assign wireOut[219] = wireIn[219];    
  assign wireOut[220] = wireIn[220];    
  assign wireOut[221] = wireIn[222];    
  assign wireOut[222] = wireIn[221];    
  assign wireOut[223] = wireIn[223];    
  assign wireOut[224] = wireIn[224];    
  assign wireOut[225] = wireIn[226];    
  assign wireOut[226] = wireIn[225];    
  assign wireOut[227] = wireIn[227];    
  assign wireOut[228] = wireIn[228];    
  assign wireOut[229] = wireIn[230];    
  assign wireOut[230] = wireIn[229];    
  assign wireOut[231] = wireIn[231];    
  assign wireOut[232] = wireIn[232];    
  assign wireOut[233] = wireIn[234];    
  assign wireOut[234] = wireIn[233];    
  assign wireOut[235] = wireIn[235];    
  assign wireOut[236] = wireIn[236];    
  assign wireOut[237] = wireIn[238];    
  assign wireOut[238] = wireIn[237];    
  assign wireOut[239] = wireIn[239];    
  assign wireOut[240] = wireIn[240];    
  assign wireOut[241] = wireIn[242];    
  assign wireOut[242] = wireIn[241];    
  assign wireOut[243] = wireIn[243];    
  assign wireOut[244] = wireIn[244];    
  assign wireOut[245] = wireIn[246];    
  assign wireOut[246] = wireIn[245];    
  assign wireOut[247] = wireIn[247];    
  assign wireOut[248] = wireIn[248];    
  assign wireOut[249] = wireIn[250];    
  assign wireOut[250] = wireIn[249];    
  assign wireOut[251] = wireIn[251];    
  assign wireOut[252] = wireIn[252];    
  assign wireOut[253] = wireIn[254];    
  assign wireOut[254] = wireIn[253];    
  assign wireOut[255] = wireIn[255];    
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module switches_stage_st7_0_L(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
ctrl,                            
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;                   
  input [128-1:0] ctrl;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  switch_2_2 switch_inst_0(.inData_0(wireIn[0]), .inData_1(wireIn[1]), .outData_0(wireOut[0]), .outData_1(wireOut[1]), .ctrl(ctrl[0]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_1(.inData_0(wireIn[2]), .inData_1(wireIn[3]), .outData_0(wireOut[2]), .outData_1(wireOut[3]), .ctrl(ctrl[1]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_2(.inData_0(wireIn[4]), .inData_1(wireIn[5]), .outData_0(wireOut[4]), .outData_1(wireOut[5]), .ctrl(ctrl[2]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_3(.inData_0(wireIn[6]), .inData_1(wireIn[7]), .outData_0(wireOut[6]), .outData_1(wireOut[7]), .ctrl(ctrl[3]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_4(.inData_0(wireIn[8]), .inData_1(wireIn[9]), .outData_0(wireOut[8]), .outData_1(wireOut[9]), .ctrl(ctrl[4]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_5(.inData_0(wireIn[10]), .inData_1(wireIn[11]), .outData_0(wireOut[10]), .outData_1(wireOut[11]), .ctrl(ctrl[5]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_6(.inData_0(wireIn[12]), .inData_1(wireIn[13]), .outData_0(wireOut[12]), .outData_1(wireOut[13]), .ctrl(ctrl[6]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_7(.inData_0(wireIn[14]), .inData_1(wireIn[15]), .outData_0(wireOut[14]), .outData_1(wireOut[15]), .ctrl(ctrl[7]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_8(.inData_0(wireIn[16]), .inData_1(wireIn[17]), .outData_0(wireOut[16]), .outData_1(wireOut[17]), .ctrl(ctrl[8]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_9(.inData_0(wireIn[18]), .inData_1(wireIn[19]), .outData_0(wireOut[18]), .outData_1(wireOut[19]), .ctrl(ctrl[9]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_10(.inData_0(wireIn[20]), .inData_1(wireIn[21]), .outData_0(wireOut[20]), .outData_1(wireOut[21]), .ctrl(ctrl[10]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_11(.inData_0(wireIn[22]), .inData_1(wireIn[23]), .outData_0(wireOut[22]), .outData_1(wireOut[23]), .ctrl(ctrl[11]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_12(.inData_0(wireIn[24]), .inData_1(wireIn[25]), .outData_0(wireOut[24]), .outData_1(wireOut[25]), .ctrl(ctrl[12]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_13(.inData_0(wireIn[26]), .inData_1(wireIn[27]), .outData_0(wireOut[26]), .outData_1(wireOut[27]), .ctrl(ctrl[13]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_14(.inData_0(wireIn[28]), .inData_1(wireIn[29]), .outData_0(wireOut[28]), .outData_1(wireOut[29]), .ctrl(ctrl[14]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_15(.inData_0(wireIn[30]), .inData_1(wireIn[31]), .outData_0(wireOut[30]), .outData_1(wireOut[31]), .ctrl(ctrl[15]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_16(.inData_0(wireIn[32]), .inData_1(wireIn[33]), .outData_0(wireOut[32]), .outData_1(wireOut[33]), .ctrl(ctrl[16]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_17(.inData_0(wireIn[34]), .inData_1(wireIn[35]), .outData_0(wireOut[34]), .outData_1(wireOut[35]), .ctrl(ctrl[17]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_18(.inData_0(wireIn[36]), .inData_1(wireIn[37]), .outData_0(wireOut[36]), .outData_1(wireOut[37]), .ctrl(ctrl[18]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_19(.inData_0(wireIn[38]), .inData_1(wireIn[39]), .outData_0(wireOut[38]), .outData_1(wireOut[39]), .ctrl(ctrl[19]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_20(.inData_0(wireIn[40]), .inData_1(wireIn[41]), .outData_0(wireOut[40]), .outData_1(wireOut[41]), .ctrl(ctrl[20]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_21(.inData_0(wireIn[42]), .inData_1(wireIn[43]), .outData_0(wireOut[42]), .outData_1(wireOut[43]), .ctrl(ctrl[21]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_22(.inData_0(wireIn[44]), .inData_1(wireIn[45]), .outData_0(wireOut[44]), .outData_1(wireOut[45]), .ctrl(ctrl[22]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_23(.inData_0(wireIn[46]), .inData_1(wireIn[47]), .outData_0(wireOut[46]), .outData_1(wireOut[47]), .ctrl(ctrl[23]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_24(.inData_0(wireIn[48]), .inData_1(wireIn[49]), .outData_0(wireOut[48]), .outData_1(wireOut[49]), .ctrl(ctrl[24]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_25(.inData_0(wireIn[50]), .inData_1(wireIn[51]), .outData_0(wireOut[50]), .outData_1(wireOut[51]), .ctrl(ctrl[25]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_26(.inData_0(wireIn[52]), .inData_1(wireIn[53]), .outData_0(wireOut[52]), .outData_1(wireOut[53]), .ctrl(ctrl[26]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_27(.inData_0(wireIn[54]), .inData_1(wireIn[55]), .outData_0(wireOut[54]), .outData_1(wireOut[55]), .ctrl(ctrl[27]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_28(.inData_0(wireIn[56]), .inData_1(wireIn[57]), .outData_0(wireOut[56]), .outData_1(wireOut[57]), .ctrl(ctrl[28]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_29(.inData_0(wireIn[58]), .inData_1(wireIn[59]), .outData_0(wireOut[58]), .outData_1(wireOut[59]), .ctrl(ctrl[29]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_30(.inData_0(wireIn[60]), .inData_1(wireIn[61]), .outData_0(wireOut[60]), .outData_1(wireOut[61]), .ctrl(ctrl[30]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_31(.inData_0(wireIn[62]), .inData_1(wireIn[63]), .outData_0(wireOut[62]), .outData_1(wireOut[63]), .ctrl(ctrl[31]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_32(.inData_0(wireIn[64]), .inData_1(wireIn[65]), .outData_0(wireOut[64]), .outData_1(wireOut[65]), .ctrl(ctrl[32]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_33(.inData_0(wireIn[66]), .inData_1(wireIn[67]), .outData_0(wireOut[66]), .outData_1(wireOut[67]), .ctrl(ctrl[33]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_34(.inData_0(wireIn[68]), .inData_1(wireIn[69]), .outData_0(wireOut[68]), .outData_1(wireOut[69]), .ctrl(ctrl[34]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_35(.inData_0(wireIn[70]), .inData_1(wireIn[71]), .outData_0(wireOut[70]), .outData_1(wireOut[71]), .ctrl(ctrl[35]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_36(.inData_0(wireIn[72]), .inData_1(wireIn[73]), .outData_0(wireOut[72]), .outData_1(wireOut[73]), .ctrl(ctrl[36]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_37(.inData_0(wireIn[74]), .inData_1(wireIn[75]), .outData_0(wireOut[74]), .outData_1(wireOut[75]), .ctrl(ctrl[37]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_38(.inData_0(wireIn[76]), .inData_1(wireIn[77]), .outData_0(wireOut[76]), .outData_1(wireOut[77]), .ctrl(ctrl[38]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_39(.inData_0(wireIn[78]), .inData_1(wireIn[79]), .outData_0(wireOut[78]), .outData_1(wireOut[79]), .ctrl(ctrl[39]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_40(.inData_0(wireIn[80]), .inData_1(wireIn[81]), .outData_0(wireOut[80]), .outData_1(wireOut[81]), .ctrl(ctrl[40]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_41(.inData_0(wireIn[82]), .inData_1(wireIn[83]), .outData_0(wireOut[82]), .outData_1(wireOut[83]), .ctrl(ctrl[41]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_42(.inData_0(wireIn[84]), .inData_1(wireIn[85]), .outData_0(wireOut[84]), .outData_1(wireOut[85]), .ctrl(ctrl[42]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_43(.inData_0(wireIn[86]), .inData_1(wireIn[87]), .outData_0(wireOut[86]), .outData_1(wireOut[87]), .ctrl(ctrl[43]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_44(.inData_0(wireIn[88]), .inData_1(wireIn[89]), .outData_0(wireOut[88]), .outData_1(wireOut[89]), .ctrl(ctrl[44]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_45(.inData_0(wireIn[90]), .inData_1(wireIn[91]), .outData_0(wireOut[90]), .outData_1(wireOut[91]), .ctrl(ctrl[45]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_46(.inData_0(wireIn[92]), .inData_1(wireIn[93]), .outData_0(wireOut[92]), .outData_1(wireOut[93]), .ctrl(ctrl[46]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_47(.inData_0(wireIn[94]), .inData_1(wireIn[95]), .outData_0(wireOut[94]), .outData_1(wireOut[95]), .ctrl(ctrl[47]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_48(.inData_0(wireIn[96]), .inData_1(wireIn[97]), .outData_0(wireOut[96]), .outData_1(wireOut[97]), .ctrl(ctrl[48]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_49(.inData_0(wireIn[98]), .inData_1(wireIn[99]), .outData_0(wireOut[98]), .outData_1(wireOut[99]), .ctrl(ctrl[49]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_50(.inData_0(wireIn[100]), .inData_1(wireIn[101]), .outData_0(wireOut[100]), .outData_1(wireOut[101]), .ctrl(ctrl[50]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_51(.inData_0(wireIn[102]), .inData_1(wireIn[103]), .outData_0(wireOut[102]), .outData_1(wireOut[103]), .ctrl(ctrl[51]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_52(.inData_0(wireIn[104]), .inData_1(wireIn[105]), .outData_0(wireOut[104]), .outData_1(wireOut[105]), .ctrl(ctrl[52]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_53(.inData_0(wireIn[106]), .inData_1(wireIn[107]), .outData_0(wireOut[106]), .outData_1(wireOut[107]), .ctrl(ctrl[53]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_54(.inData_0(wireIn[108]), .inData_1(wireIn[109]), .outData_0(wireOut[108]), .outData_1(wireOut[109]), .ctrl(ctrl[54]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_55(.inData_0(wireIn[110]), .inData_1(wireIn[111]), .outData_0(wireOut[110]), .outData_1(wireOut[111]), .ctrl(ctrl[55]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_56(.inData_0(wireIn[112]), .inData_1(wireIn[113]), .outData_0(wireOut[112]), .outData_1(wireOut[113]), .ctrl(ctrl[56]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_57(.inData_0(wireIn[114]), .inData_1(wireIn[115]), .outData_0(wireOut[114]), .outData_1(wireOut[115]), .ctrl(ctrl[57]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_58(.inData_0(wireIn[116]), .inData_1(wireIn[117]), .outData_0(wireOut[116]), .outData_1(wireOut[117]), .ctrl(ctrl[58]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_59(.inData_0(wireIn[118]), .inData_1(wireIn[119]), .outData_0(wireOut[118]), .outData_1(wireOut[119]), .ctrl(ctrl[59]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_60(.inData_0(wireIn[120]), .inData_1(wireIn[121]), .outData_0(wireOut[120]), .outData_1(wireOut[121]), .ctrl(ctrl[60]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_61(.inData_0(wireIn[122]), .inData_1(wireIn[123]), .outData_0(wireOut[122]), .outData_1(wireOut[123]), .ctrl(ctrl[61]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_62(.inData_0(wireIn[124]), .inData_1(wireIn[125]), .outData_0(wireOut[124]), .outData_1(wireOut[125]), .ctrl(ctrl[62]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_63(.inData_0(wireIn[126]), .inData_1(wireIn[127]), .outData_0(wireOut[126]), .outData_1(wireOut[127]), .ctrl(ctrl[63]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_64(.inData_0(wireIn[128]), .inData_1(wireIn[129]), .outData_0(wireOut[128]), .outData_1(wireOut[129]), .ctrl(ctrl[64]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_65(.inData_0(wireIn[130]), .inData_1(wireIn[131]), .outData_0(wireOut[130]), .outData_1(wireOut[131]), .ctrl(ctrl[65]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_66(.inData_0(wireIn[132]), .inData_1(wireIn[133]), .outData_0(wireOut[132]), .outData_1(wireOut[133]), .ctrl(ctrl[66]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_67(.inData_0(wireIn[134]), .inData_1(wireIn[135]), .outData_0(wireOut[134]), .outData_1(wireOut[135]), .ctrl(ctrl[67]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_68(.inData_0(wireIn[136]), .inData_1(wireIn[137]), .outData_0(wireOut[136]), .outData_1(wireOut[137]), .ctrl(ctrl[68]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_69(.inData_0(wireIn[138]), .inData_1(wireIn[139]), .outData_0(wireOut[138]), .outData_1(wireOut[139]), .ctrl(ctrl[69]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_70(.inData_0(wireIn[140]), .inData_1(wireIn[141]), .outData_0(wireOut[140]), .outData_1(wireOut[141]), .ctrl(ctrl[70]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_71(.inData_0(wireIn[142]), .inData_1(wireIn[143]), .outData_0(wireOut[142]), .outData_1(wireOut[143]), .ctrl(ctrl[71]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_72(.inData_0(wireIn[144]), .inData_1(wireIn[145]), .outData_0(wireOut[144]), .outData_1(wireOut[145]), .ctrl(ctrl[72]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_73(.inData_0(wireIn[146]), .inData_1(wireIn[147]), .outData_0(wireOut[146]), .outData_1(wireOut[147]), .ctrl(ctrl[73]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_74(.inData_0(wireIn[148]), .inData_1(wireIn[149]), .outData_0(wireOut[148]), .outData_1(wireOut[149]), .ctrl(ctrl[74]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_75(.inData_0(wireIn[150]), .inData_1(wireIn[151]), .outData_0(wireOut[150]), .outData_1(wireOut[151]), .ctrl(ctrl[75]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_76(.inData_0(wireIn[152]), .inData_1(wireIn[153]), .outData_0(wireOut[152]), .outData_1(wireOut[153]), .ctrl(ctrl[76]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_77(.inData_0(wireIn[154]), .inData_1(wireIn[155]), .outData_0(wireOut[154]), .outData_1(wireOut[155]), .ctrl(ctrl[77]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_78(.inData_0(wireIn[156]), .inData_1(wireIn[157]), .outData_0(wireOut[156]), .outData_1(wireOut[157]), .ctrl(ctrl[78]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_79(.inData_0(wireIn[158]), .inData_1(wireIn[159]), .outData_0(wireOut[158]), .outData_1(wireOut[159]), .ctrl(ctrl[79]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_80(.inData_0(wireIn[160]), .inData_1(wireIn[161]), .outData_0(wireOut[160]), .outData_1(wireOut[161]), .ctrl(ctrl[80]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_81(.inData_0(wireIn[162]), .inData_1(wireIn[163]), .outData_0(wireOut[162]), .outData_1(wireOut[163]), .ctrl(ctrl[81]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_82(.inData_0(wireIn[164]), .inData_1(wireIn[165]), .outData_0(wireOut[164]), .outData_1(wireOut[165]), .ctrl(ctrl[82]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_83(.inData_0(wireIn[166]), .inData_1(wireIn[167]), .outData_0(wireOut[166]), .outData_1(wireOut[167]), .ctrl(ctrl[83]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_84(.inData_0(wireIn[168]), .inData_1(wireIn[169]), .outData_0(wireOut[168]), .outData_1(wireOut[169]), .ctrl(ctrl[84]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_85(.inData_0(wireIn[170]), .inData_1(wireIn[171]), .outData_0(wireOut[170]), .outData_1(wireOut[171]), .ctrl(ctrl[85]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_86(.inData_0(wireIn[172]), .inData_1(wireIn[173]), .outData_0(wireOut[172]), .outData_1(wireOut[173]), .ctrl(ctrl[86]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_87(.inData_0(wireIn[174]), .inData_1(wireIn[175]), .outData_0(wireOut[174]), .outData_1(wireOut[175]), .ctrl(ctrl[87]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_88(.inData_0(wireIn[176]), .inData_1(wireIn[177]), .outData_0(wireOut[176]), .outData_1(wireOut[177]), .ctrl(ctrl[88]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_89(.inData_0(wireIn[178]), .inData_1(wireIn[179]), .outData_0(wireOut[178]), .outData_1(wireOut[179]), .ctrl(ctrl[89]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_90(.inData_0(wireIn[180]), .inData_1(wireIn[181]), .outData_0(wireOut[180]), .outData_1(wireOut[181]), .ctrl(ctrl[90]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_91(.inData_0(wireIn[182]), .inData_1(wireIn[183]), .outData_0(wireOut[182]), .outData_1(wireOut[183]), .ctrl(ctrl[91]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_92(.inData_0(wireIn[184]), .inData_1(wireIn[185]), .outData_0(wireOut[184]), .outData_1(wireOut[185]), .ctrl(ctrl[92]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_93(.inData_0(wireIn[186]), .inData_1(wireIn[187]), .outData_0(wireOut[186]), .outData_1(wireOut[187]), .ctrl(ctrl[93]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_94(.inData_0(wireIn[188]), .inData_1(wireIn[189]), .outData_0(wireOut[188]), .outData_1(wireOut[189]), .ctrl(ctrl[94]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_95(.inData_0(wireIn[190]), .inData_1(wireIn[191]), .outData_0(wireOut[190]), .outData_1(wireOut[191]), .ctrl(ctrl[95]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_96(.inData_0(wireIn[192]), .inData_1(wireIn[193]), .outData_0(wireOut[192]), .outData_1(wireOut[193]), .ctrl(ctrl[96]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_97(.inData_0(wireIn[194]), .inData_1(wireIn[195]), .outData_0(wireOut[194]), .outData_1(wireOut[195]), .ctrl(ctrl[97]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_98(.inData_0(wireIn[196]), .inData_1(wireIn[197]), .outData_0(wireOut[196]), .outData_1(wireOut[197]), .ctrl(ctrl[98]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_99(.inData_0(wireIn[198]), .inData_1(wireIn[199]), .outData_0(wireOut[198]), .outData_1(wireOut[199]), .ctrl(ctrl[99]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_100(.inData_0(wireIn[200]), .inData_1(wireIn[201]), .outData_0(wireOut[200]), .outData_1(wireOut[201]), .ctrl(ctrl[100]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_101(.inData_0(wireIn[202]), .inData_1(wireIn[203]), .outData_0(wireOut[202]), .outData_1(wireOut[203]), .ctrl(ctrl[101]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_102(.inData_0(wireIn[204]), .inData_1(wireIn[205]), .outData_0(wireOut[204]), .outData_1(wireOut[205]), .ctrl(ctrl[102]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_103(.inData_0(wireIn[206]), .inData_1(wireIn[207]), .outData_0(wireOut[206]), .outData_1(wireOut[207]), .ctrl(ctrl[103]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_104(.inData_0(wireIn[208]), .inData_1(wireIn[209]), .outData_0(wireOut[208]), .outData_1(wireOut[209]), .ctrl(ctrl[104]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_105(.inData_0(wireIn[210]), .inData_1(wireIn[211]), .outData_0(wireOut[210]), .outData_1(wireOut[211]), .ctrl(ctrl[105]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_106(.inData_0(wireIn[212]), .inData_1(wireIn[213]), .outData_0(wireOut[212]), .outData_1(wireOut[213]), .ctrl(ctrl[106]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_107(.inData_0(wireIn[214]), .inData_1(wireIn[215]), .outData_0(wireOut[214]), .outData_1(wireOut[215]), .ctrl(ctrl[107]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_108(.inData_0(wireIn[216]), .inData_1(wireIn[217]), .outData_0(wireOut[216]), .outData_1(wireOut[217]), .ctrl(ctrl[108]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_109(.inData_0(wireIn[218]), .inData_1(wireIn[219]), .outData_0(wireOut[218]), .outData_1(wireOut[219]), .ctrl(ctrl[109]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_110(.inData_0(wireIn[220]), .inData_1(wireIn[221]), .outData_0(wireOut[220]), .outData_1(wireOut[221]), .ctrl(ctrl[110]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_111(.inData_0(wireIn[222]), .inData_1(wireIn[223]), .outData_0(wireOut[222]), .outData_1(wireOut[223]), .ctrl(ctrl[111]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_112(.inData_0(wireIn[224]), .inData_1(wireIn[225]), .outData_0(wireOut[224]), .outData_1(wireOut[225]), .ctrl(ctrl[112]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_113(.inData_0(wireIn[226]), .inData_1(wireIn[227]), .outData_0(wireOut[226]), .outData_1(wireOut[227]), .ctrl(ctrl[113]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_114(.inData_0(wireIn[228]), .inData_1(wireIn[229]), .outData_0(wireOut[228]), .outData_1(wireOut[229]), .ctrl(ctrl[114]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_115(.inData_0(wireIn[230]), .inData_1(wireIn[231]), .outData_0(wireOut[230]), .outData_1(wireOut[231]), .ctrl(ctrl[115]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_116(.inData_0(wireIn[232]), .inData_1(wireIn[233]), .outData_0(wireOut[232]), .outData_1(wireOut[233]), .ctrl(ctrl[116]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_117(.inData_0(wireIn[234]), .inData_1(wireIn[235]), .outData_0(wireOut[234]), .outData_1(wireOut[235]), .ctrl(ctrl[117]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_118(.inData_0(wireIn[236]), .inData_1(wireIn[237]), .outData_0(wireOut[236]), .outData_1(wireOut[237]), .ctrl(ctrl[118]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_119(.inData_0(wireIn[238]), .inData_1(wireIn[239]), .outData_0(wireOut[238]), .outData_1(wireOut[239]), .ctrl(ctrl[119]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_120(.inData_0(wireIn[240]), .inData_1(wireIn[241]), .outData_0(wireOut[240]), .outData_1(wireOut[241]), .ctrl(ctrl[120]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_121(.inData_0(wireIn[242]), .inData_1(wireIn[243]), .outData_0(wireOut[242]), .outData_1(wireOut[243]), .ctrl(ctrl[121]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_122(.inData_0(wireIn[244]), .inData_1(wireIn[245]), .outData_0(wireOut[244]), .outData_1(wireOut[245]), .ctrl(ctrl[122]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_123(.inData_0(wireIn[246]), .inData_1(wireIn[247]), .outData_0(wireOut[246]), .outData_1(wireOut[247]), .ctrl(ctrl[123]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_124(.inData_0(wireIn[248]), .inData_1(wireIn[249]), .outData_0(wireOut[248]), .outData_1(wireOut[249]), .ctrl(ctrl[124]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_125(.inData_0(wireIn[250]), .inData_1(wireIn[251]), .outData_0(wireOut[250]), .outData_1(wireOut[251]), .ctrl(ctrl[125]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_126(.inData_0(wireIn[252]), .inData_1(wireIn[253]), .outData_0(wireOut[252]), .outData_1(wireOut[253]), .ctrl(ctrl[126]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_127(.inData_0(wireIn[254]), .inData_1(wireIn[255]), .outData_0(wireOut[254]), .outData_1(wireOut[255]), .ctrl(ctrl[127]), .clk(clk), .rst(rst));
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module wireCon_dp256_st7_L(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  assign wireOut[0] = wireIn[0];    
  assign wireOut[1] = wireIn[1];    
  assign wireOut[2] = wireIn[2];    
  assign wireOut[3] = wireIn[3];    
  assign wireOut[4] = wireIn[4];    
  assign wireOut[5] = wireIn[5];    
  assign wireOut[6] = wireIn[6];    
  assign wireOut[7] = wireIn[7];    
  assign wireOut[8] = wireIn[8];    
  assign wireOut[9] = wireIn[9];    
  assign wireOut[10] = wireIn[10];    
  assign wireOut[11] = wireIn[11];    
  assign wireOut[12] = wireIn[12];    
  assign wireOut[13] = wireIn[13];    
  assign wireOut[14] = wireIn[14];    
  assign wireOut[15] = wireIn[15];    
  assign wireOut[16] = wireIn[16];    
  assign wireOut[17] = wireIn[17];    
  assign wireOut[18] = wireIn[18];    
  assign wireOut[19] = wireIn[19];    
  assign wireOut[20] = wireIn[20];    
  assign wireOut[21] = wireIn[21];    
  assign wireOut[22] = wireIn[22];    
  assign wireOut[23] = wireIn[23];    
  assign wireOut[24] = wireIn[24];    
  assign wireOut[25] = wireIn[25];    
  assign wireOut[26] = wireIn[26];    
  assign wireOut[27] = wireIn[27];    
  assign wireOut[28] = wireIn[28];    
  assign wireOut[29] = wireIn[29];    
  assign wireOut[30] = wireIn[30];    
  assign wireOut[31] = wireIn[31];    
  assign wireOut[32] = wireIn[32];    
  assign wireOut[33] = wireIn[33];    
  assign wireOut[34] = wireIn[34];    
  assign wireOut[35] = wireIn[35];    
  assign wireOut[36] = wireIn[36];    
  assign wireOut[37] = wireIn[37];    
  assign wireOut[38] = wireIn[38];    
  assign wireOut[39] = wireIn[39];    
  assign wireOut[40] = wireIn[40];    
  assign wireOut[41] = wireIn[41];    
  assign wireOut[42] = wireIn[42];    
  assign wireOut[43] = wireIn[43];    
  assign wireOut[44] = wireIn[44];    
  assign wireOut[45] = wireIn[45];    
  assign wireOut[46] = wireIn[46];    
  assign wireOut[47] = wireIn[47];    
  assign wireOut[48] = wireIn[48];    
  assign wireOut[49] = wireIn[49];    
  assign wireOut[50] = wireIn[50];    
  assign wireOut[51] = wireIn[51];    
  assign wireOut[52] = wireIn[52];    
  assign wireOut[53] = wireIn[53];    
  assign wireOut[54] = wireIn[54];    
  assign wireOut[55] = wireIn[55];    
  assign wireOut[56] = wireIn[56];    
  assign wireOut[57] = wireIn[57];    
  assign wireOut[58] = wireIn[58];    
  assign wireOut[59] = wireIn[59];    
  assign wireOut[60] = wireIn[60];    
  assign wireOut[61] = wireIn[61];    
  assign wireOut[62] = wireIn[62];    
  assign wireOut[63] = wireIn[63];    
  assign wireOut[64] = wireIn[64];    
  assign wireOut[65] = wireIn[65];    
  assign wireOut[66] = wireIn[66];    
  assign wireOut[67] = wireIn[67];    
  assign wireOut[68] = wireIn[68];    
  assign wireOut[69] = wireIn[69];    
  assign wireOut[70] = wireIn[70];    
  assign wireOut[71] = wireIn[71];    
  assign wireOut[72] = wireIn[72];    
  assign wireOut[73] = wireIn[73];    
  assign wireOut[74] = wireIn[74];    
  assign wireOut[75] = wireIn[75];    
  assign wireOut[76] = wireIn[76];    
  assign wireOut[77] = wireIn[77];    
  assign wireOut[78] = wireIn[78];    
  assign wireOut[79] = wireIn[79];    
  assign wireOut[80] = wireIn[80];    
  assign wireOut[81] = wireIn[81];    
  assign wireOut[82] = wireIn[82];    
  assign wireOut[83] = wireIn[83];    
  assign wireOut[84] = wireIn[84];    
  assign wireOut[85] = wireIn[85];    
  assign wireOut[86] = wireIn[86];    
  assign wireOut[87] = wireIn[87];    
  assign wireOut[88] = wireIn[88];    
  assign wireOut[89] = wireIn[89];    
  assign wireOut[90] = wireIn[90];    
  assign wireOut[91] = wireIn[91];    
  assign wireOut[92] = wireIn[92];    
  assign wireOut[93] = wireIn[93];    
  assign wireOut[94] = wireIn[94];    
  assign wireOut[95] = wireIn[95];    
  assign wireOut[96] = wireIn[96];    
  assign wireOut[97] = wireIn[97];    
  assign wireOut[98] = wireIn[98];    
  assign wireOut[99] = wireIn[99];    
  assign wireOut[100] = wireIn[100];    
  assign wireOut[101] = wireIn[101];    
  assign wireOut[102] = wireIn[102];    
  assign wireOut[103] = wireIn[103];    
  assign wireOut[104] = wireIn[104];    
  assign wireOut[105] = wireIn[105];    
  assign wireOut[106] = wireIn[106];    
  assign wireOut[107] = wireIn[107];    
  assign wireOut[108] = wireIn[108];    
  assign wireOut[109] = wireIn[109];    
  assign wireOut[110] = wireIn[110];    
  assign wireOut[111] = wireIn[111];    
  assign wireOut[112] = wireIn[112];    
  assign wireOut[113] = wireIn[113];    
  assign wireOut[114] = wireIn[114];    
  assign wireOut[115] = wireIn[115];    
  assign wireOut[116] = wireIn[116];    
  assign wireOut[117] = wireIn[117];    
  assign wireOut[118] = wireIn[118];    
  assign wireOut[119] = wireIn[119];    
  assign wireOut[120] = wireIn[120];    
  assign wireOut[121] = wireIn[121];    
  assign wireOut[122] = wireIn[122];    
  assign wireOut[123] = wireIn[123];    
  assign wireOut[124] = wireIn[124];    
  assign wireOut[125] = wireIn[125];    
  assign wireOut[126] = wireIn[126];    
  assign wireOut[127] = wireIn[127];    
  assign wireOut[128] = wireIn[128];    
  assign wireOut[129] = wireIn[129];    
  assign wireOut[130] = wireIn[130];    
  assign wireOut[131] = wireIn[131];    
  assign wireOut[132] = wireIn[132];    
  assign wireOut[133] = wireIn[133];    
  assign wireOut[134] = wireIn[134];    
  assign wireOut[135] = wireIn[135];    
  assign wireOut[136] = wireIn[136];    
  assign wireOut[137] = wireIn[137];    
  assign wireOut[138] = wireIn[138];    
  assign wireOut[139] = wireIn[139];    
  assign wireOut[140] = wireIn[140];    
  assign wireOut[141] = wireIn[141];    
  assign wireOut[142] = wireIn[142];    
  assign wireOut[143] = wireIn[143];    
  assign wireOut[144] = wireIn[144];    
  assign wireOut[145] = wireIn[145];    
  assign wireOut[146] = wireIn[146];    
  assign wireOut[147] = wireIn[147];    
  assign wireOut[148] = wireIn[148];    
  assign wireOut[149] = wireIn[149];    
  assign wireOut[150] = wireIn[150];    
  assign wireOut[151] = wireIn[151];    
  assign wireOut[152] = wireIn[152];    
  assign wireOut[153] = wireIn[153];    
  assign wireOut[154] = wireIn[154];    
  assign wireOut[155] = wireIn[155];    
  assign wireOut[156] = wireIn[156];    
  assign wireOut[157] = wireIn[157];    
  assign wireOut[158] = wireIn[158];    
  assign wireOut[159] = wireIn[159];    
  assign wireOut[160] = wireIn[160];    
  assign wireOut[161] = wireIn[161];    
  assign wireOut[162] = wireIn[162];    
  assign wireOut[163] = wireIn[163];    
  assign wireOut[164] = wireIn[164];    
  assign wireOut[165] = wireIn[165];    
  assign wireOut[166] = wireIn[166];    
  assign wireOut[167] = wireIn[167];    
  assign wireOut[168] = wireIn[168];    
  assign wireOut[169] = wireIn[169];    
  assign wireOut[170] = wireIn[170];    
  assign wireOut[171] = wireIn[171];    
  assign wireOut[172] = wireIn[172];    
  assign wireOut[173] = wireIn[173];    
  assign wireOut[174] = wireIn[174];    
  assign wireOut[175] = wireIn[175];    
  assign wireOut[176] = wireIn[176];    
  assign wireOut[177] = wireIn[177];    
  assign wireOut[178] = wireIn[178];    
  assign wireOut[179] = wireIn[179];    
  assign wireOut[180] = wireIn[180];    
  assign wireOut[181] = wireIn[181];    
  assign wireOut[182] = wireIn[182];    
  assign wireOut[183] = wireIn[183];    
  assign wireOut[184] = wireIn[184];    
  assign wireOut[185] = wireIn[185];    
  assign wireOut[186] = wireIn[186];    
  assign wireOut[187] = wireIn[187];    
  assign wireOut[188] = wireIn[188];    
  assign wireOut[189] = wireIn[189];    
  assign wireOut[190] = wireIn[190];    
  assign wireOut[191] = wireIn[191];    
  assign wireOut[192] = wireIn[192];    
  assign wireOut[193] = wireIn[193];    
  assign wireOut[194] = wireIn[194];    
  assign wireOut[195] = wireIn[195];    
  assign wireOut[196] = wireIn[196];    
  assign wireOut[197] = wireIn[197];    
  assign wireOut[198] = wireIn[198];    
  assign wireOut[199] = wireIn[199];    
  assign wireOut[200] = wireIn[200];    
  assign wireOut[201] = wireIn[201];    
  assign wireOut[202] = wireIn[202];    
  assign wireOut[203] = wireIn[203];    
  assign wireOut[204] = wireIn[204];    
  assign wireOut[205] = wireIn[205];    
  assign wireOut[206] = wireIn[206];    
  assign wireOut[207] = wireIn[207];    
  assign wireOut[208] = wireIn[208];    
  assign wireOut[209] = wireIn[209];    
  assign wireOut[210] = wireIn[210];    
  assign wireOut[211] = wireIn[211];    
  assign wireOut[212] = wireIn[212];    
  assign wireOut[213] = wireIn[213];    
  assign wireOut[214] = wireIn[214];    
  assign wireOut[215] = wireIn[215];    
  assign wireOut[216] = wireIn[216];    
  assign wireOut[217] = wireIn[217];    
  assign wireOut[218] = wireIn[218];    
  assign wireOut[219] = wireIn[219];    
  assign wireOut[220] = wireIn[220];    
  assign wireOut[221] = wireIn[221];    
  assign wireOut[222] = wireIn[222];    
  assign wireOut[223] = wireIn[223];    
  assign wireOut[224] = wireIn[224];    
  assign wireOut[225] = wireIn[225];    
  assign wireOut[226] = wireIn[226];    
  assign wireOut[227] = wireIn[227];    
  assign wireOut[228] = wireIn[228];    
  assign wireOut[229] = wireIn[229];    
  assign wireOut[230] = wireIn[230];    
  assign wireOut[231] = wireIn[231];    
  assign wireOut[232] = wireIn[232];    
  assign wireOut[233] = wireIn[233];    
  assign wireOut[234] = wireIn[234];    
  assign wireOut[235] = wireIn[235];    
  assign wireOut[236] = wireIn[236];    
  assign wireOut[237] = wireIn[237];    
  assign wireOut[238] = wireIn[238];    
  assign wireOut[239] = wireIn[239];    
  assign wireOut[240] = wireIn[240];    
  assign wireOut[241] = wireIn[241];    
  assign wireOut[242] = wireIn[242];    
  assign wireOut[243] = wireIn[243];    
  assign wireOut[244] = wireIn[244];    
  assign wireOut[245] = wireIn[245];    
  assign wireOut[246] = wireIn[246];    
  assign wireOut[247] = wireIn[247];    
  assign wireOut[248] = wireIn[248];    
  assign wireOut[249] = wireIn[249];    
  assign wireOut[250] = wireIn[250];    
  assign wireOut[251] = wireIn[251];    
  assign wireOut[252] = wireIn[252];    
  assign wireOut[253] = wireIn[253];    
  assign wireOut[254] = wireIn[254];    
  assign wireOut[255] = wireIn[255];    
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module ingressStage_p256(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
counter_in,                       
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;                   
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  input [7:0] counter_in; 
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255;
  output out_start; 
  
  
  wire out_start_w; 
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  wire in_start_stage0;
  wire con_in_start_stage0;

  wire in_start_stage1;
  wire con_in_start_stage1;

  wire in_start_stage2;
  wire con_in_start_stage2;

  wire in_start_stage3;
  wire con_in_start_stage3;

  wire in_start_stage4;
  wire con_in_start_stage4;

  wire in_start_stage5;
  wire con_in_start_stage5;

  wire in_start_stage6;
  wire con_in_start_stage6;

  wire in_start_stage7;
  wire con_in_start_stage7;

  wire [DATA_WIDTH-1:0] wire_con_in_stage0[255:0];
  wire [DATA_WIDTH-1:0] wire_con_out_stage0[255:0];
  wire [127:0] wire_ctrl_stage0;

  switches_stage_st0_0_L switch_stage_0(
        .inData_0(wireIn[0]), .inData_1(wireIn[1]), .inData_2(wireIn[2]), .inData_3(wireIn[3]), .inData_4(wireIn[4]), .inData_5(wireIn[5]), .inData_6(wireIn[6]), .inData_7(wireIn[7]), .inData_8(wireIn[8]), .inData_9(wireIn[9]), .inData_10(wireIn[10]), .inData_11(wireIn[11]), .inData_12(wireIn[12]), .inData_13(wireIn[13]), .inData_14(wireIn[14]), .inData_15(wireIn[15]), .inData_16(wireIn[16]), .inData_17(wireIn[17]), .inData_18(wireIn[18]), .inData_19(wireIn[19]), .inData_20(wireIn[20]), .inData_21(wireIn[21]), .inData_22(wireIn[22]), .inData_23(wireIn[23]), .inData_24(wireIn[24]), .inData_25(wireIn[25]), .inData_26(wireIn[26]), .inData_27(wireIn[27]), .inData_28(wireIn[28]), .inData_29(wireIn[29]), .inData_30(wireIn[30]), .inData_31(wireIn[31]), .inData_32(wireIn[32]), .inData_33(wireIn[33]), .inData_34(wireIn[34]), .inData_35(wireIn[35]), .inData_36(wireIn[36]), .inData_37(wireIn[37]), .inData_38(wireIn[38]), .inData_39(wireIn[39]), .inData_40(wireIn[40]), .inData_41(wireIn[41]), .inData_42(wireIn[42]), .inData_43(wireIn[43]), .inData_44(wireIn[44]), .inData_45(wireIn[45]), .inData_46(wireIn[46]), .inData_47(wireIn[47]), .inData_48(wireIn[48]), .inData_49(wireIn[49]), .inData_50(wireIn[50]), .inData_51(wireIn[51]), .inData_52(wireIn[52]), .inData_53(wireIn[53]), .inData_54(wireIn[54]), .inData_55(wireIn[55]), .inData_56(wireIn[56]), .inData_57(wireIn[57]), .inData_58(wireIn[58]), .inData_59(wireIn[59]), .inData_60(wireIn[60]), .inData_61(wireIn[61]), .inData_62(wireIn[62]), .inData_63(wireIn[63]), .inData_64(wireIn[64]), .inData_65(wireIn[65]), .inData_66(wireIn[66]), .inData_67(wireIn[67]), .inData_68(wireIn[68]), .inData_69(wireIn[69]), .inData_70(wireIn[70]), .inData_71(wireIn[71]), .inData_72(wireIn[72]), .inData_73(wireIn[73]), .inData_74(wireIn[74]), .inData_75(wireIn[75]), .inData_76(wireIn[76]), .inData_77(wireIn[77]), .inData_78(wireIn[78]), .inData_79(wireIn[79]), .inData_80(wireIn[80]), .inData_81(wireIn[81]), .inData_82(wireIn[82]), .inData_83(wireIn[83]), .inData_84(wireIn[84]), .inData_85(wireIn[85]), .inData_86(wireIn[86]), .inData_87(wireIn[87]), .inData_88(wireIn[88]), .inData_89(wireIn[89]), .inData_90(wireIn[90]), .inData_91(wireIn[91]), .inData_92(wireIn[92]), .inData_93(wireIn[93]), .inData_94(wireIn[94]), .inData_95(wireIn[95]), .inData_96(wireIn[96]), .inData_97(wireIn[97]), .inData_98(wireIn[98]), .inData_99(wireIn[99]), .inData_100(wireIn[100]), .inData_101(wireIn[101]), .inData_102(wireIn[102]), .inData_103(wireIn[103]), .inData_104(wireIn[104]), .inData_105(wireIn[105]), .inData_106(wireIn[106]), .inData_107(wireIn[107]), .inData_108(wireIn[108]), .inData_109(wireIn[109]), .inData_110(wireIn[110]), .inData_111(wireIn[111]), .inData_112(wireIn[112]), .inData_113(wireIn[113]), .inData_114(wireIn[114]), .inData_115(wireIn[115]), .inData_116(wireIn[116]), .inData_117(wireIn[117]), .inData_118(wireIn[118]), .inData_119(wireIn[119]), .inData_120(wireIn[120]), .inData_121(wireIn[121]), .inData_122(wireIn[122]), .inData_123(wireIn[123]), .inData_124(wireIn[124]), .inData_125(wireIn[125]), .inData_126(wireIn[126]), .inData_127(wireIn[127]), .inData_128(wireIn[128]), .inData_129(wireIn[129]), .inData_130(wireIn[130]), .inData_131(wireIn[131]), .inData_132(wireIn[132]), .inData_133(wireIn[133]), .inData_134(wireIn[134]), .inData_135(wireIn[135]), .inData_136(wireIn[136]), .inData_137(wireIn[137]), .inData_138(wireIn[138]), .inData_139(wireIn[139]), .inData_140(wireIn[140]), .inData_141(wireIn[141]), .inData_142(wireIn[142]), .inData_143(wireIn[143]), .inData_144(wireIn[144]), .inData_145(wireIn[145]), .inData_146(wireIn[146]), .inData_147(wireIn[147]), .inData_148(wireIn[148]), .inData_149(wireIn[149]), .inData_150(wireIn[150]), .inData_151(wireIn[151]), .inData_152(wireIn[152]), .inData_153(wireIn[153]), .inData_154(wireIn[154]), .inData_155(wireIn[155]), .inData_156(wireIn[156]), .inData_157(wireIn[157]), .inData_158(wireIn[158]), .inData_159(wireIn[159]), .inData_160(wireIn[160]), .inData_161(wireIn[161]), .inData_162(wireIn[162]), .inData_163(wireIn[163]), .inData_164(wireIn[164]), .inData_165(wireIn[165]), .inData_166(wireIn[166]), .inData_167(wireIn[167]), .inData_168(wireIn[168]), .inData_169(wireIn[169]), .inData_170(wireIn[170]), .inData_171(wireIn[171]), .inData_172(wireIn[172]), .inData_173(wireIn[173]), .inData_174(wireIn[174]), .inData_175(wireIn[175]), .inData_176(wireIn[176]), .inData_177(wireIn[177]), .inData_178(wireIn[178]), .inData_179(wireIn[179]), .inData_180(wireIn[180]), .inData_181(wireIn[181]), .inData_182(wireIn[182]), .inData_183(wireIn[183]), .inData_184(wireIn[184]), .inData_185(wireIn[185]), .inData_186(wireIn[186]), .inData_187(wireIn[187]), .inData_188(wireIn[188]), .inData_189(wireIn[189]), .inData_190(wireIn[190]), .inData_191(wireIn[191]), .inData_192(wireIn[192]), .inData_193(wireIn[193]), .inData_194(wireIn[194]), .inData_195(wireIn[195]), .inData_196(wireIn[196]), .inData_197(wireIn[197]), .inData_198(wireIn[198]), .inData_199(wireIn[199]), .inData_200(wireIn[200]), .inData_201(wireIn[201]), .inData_202(wireIn[202]), .inData_203(wireIn[203]), .inData_204(wireIn[204]), .inData_205(wireIn[205]), .inData_206(wireIn[206]), .inData_207(wireIn[207]), .inData_208(wireIn[208]), .inData_209(wireIn[209]), .inData_210(wireIn[210]), .inData_211(wireIn[211]), .inData_212(wireIn[212]), .inData_213(wireIn[213]), .inData_214(wireIn[214]), .inData_215(wireIn[215]), .inData_216(wireIn[216]), .inData_217(wireIn[217]), .inData_218(wireIn[218]), .inData_219(wireIn[219]), .inData_220(wireIn[220]), .inData_221(wireIn[221]), .inData_222(wireIn[222]), .inData_223(wireIn[223]), .inData_224(wireIn[224]), .inData_225(wireIn[225]), .inData_226(wireIn[226]), .inData_227(wireIn[227]), .inData_228(wireIn[228]), .inData_229(wireIn[229]), .inData_230(wireIn[230]), .inData_231(wireIn[231]), .inData_232(wireIn[232]), .inData_233(wireIn[233]), .inData_234(wireIn[234]), .inData_235(wireIn[235]), .inData_236(wireIn[236]), .inData_237(wireIn[237]), .inData_238(wireIn[238]), .inData_239(wireIn[239]), .inData_240(wireIn[240]), .inData_241(wireIn[241]), .inData_242(wireIn[242]), .inData_243(wireIn[243]), .inData_244(wireIn[244]), .inData_245(wireIn[245]), .inData_246(wireIn[246]), .inData_247(wireIn[247]), .inData_248(wireIn[248]), .inData_249(wireIn[249]), .inData_250(wireIn[250]), .inData_251(wireIn[251]), .inData_252(wireIn[252]), .inData_253(wireIn[253]), .inData_254(wireIn[254]), .inData_255(wireIn[255]), 
        .outData_0(wire_con_in_stage0[0]), .outData_1(wire_con_in_stage0[1]), .outData_2(wire_con_in_stage0[2]), .outData_3(wire_con_in_stage0[3]), .outData_4(wire_con_in_stage0[4]), .outData_5(wire_con_in_stage0[5]), .outData_6(wire_con_in_stage0[6]), .outData_7(wire_con_in_stage0[7]), .outData_8(wire_con_in_stage0[8]), .outData_9(wire_con_in_stage0[9]), .outData_10(wire_con_in_stage0[10]), .outData_11(wire_con_in_stage0[11]), .outData_12(wire_con_in_stage0[12]), .outData_13(wire_con_in_stage0[13]), .outData_14(wire_con_in_stage0[14]), .outData_15(wire_con_in_stage0[15]), .outData_16(wire_con_in_stage0[16]), .outData_17(wire_con_in_stage0[17]), .outData_18(wire_con_in_stage0[18]), .outData_19(wire_con_in_stage0[19]), .outData_20(wire_con_in_stage0[20]), .outData_21(wire_con_in_stage0[21]), .outData_22(wire_con_in_stage0[22]), .outData_23(wire_con_in_stage0[23]), .outData_24(wire_con_in_stage0[24]), .outData_25(wire_con_in_stage0[25]), .outData_26(wire_con_in_stage0[26]), .outData_27(wire_con_in_stage0[27]), .outData_28(wire_con_in_stage0[28]), .outData_29(wire_con_in_stage0[29]), .outData_30(wire_con_in_stage0[30]), .outData_31(wire_con_in_stage0[31]), .outData_32(wire_con_in_stage0[32]), .outData_33(wire_con_in_stage0[33]), .outData_34(wire_con_in_stage0[34]), .outData_35(wire_con_in_stage0[35]), .outData_36(wire_con_in_stage0[36]), .outData_37(wire_con_in_stage0[37]), .outData_38(wire_con_in_stage0[38]), .outData_39(wire_con_in_stage0[39]), .outData_40(wire_con_in_stage0[40]), .outData_41(wire_con_in_stage0[41]), .outData_42(wire_con_in_stage0[42]), .outData_43(wire_con_in_stage0[43]), .outData_44(wire_con_in_stage0[44]), .outData_45(wire_con_in_stage0[45]), .outData_46(wire_con_in_stage0[46]), .outData_47(wire_con_in_stage0[47]), .outData_48(wire_con_in_stage0[48]), .outData_49(wire_con_in_stage0[49]), .outData_50(wire_con_in_stage0[50]), .outData_51(wire_con_in_stage0[51]), .outData_52(wire_con_in_stage0[52]), .outData_53(wire_con_in_stage0[53]), .outData_54(wire_con_in_stage0[54]), .outData_55(wire_con_in_stage0[55]), .outData_56(wire_con_in_stage0[56]), .outData_57(wire_con_in_stage0[57]), .outData_58(wire_con_in_stage0[58]), .outData_59(wire_con_in_stage0[59]), .outData_60(wire_con_in_stage0[60]), .outData_61(wire_con_in_stage0[61]), .outData_62(wire_con_in_stage0[62]), .outData_63(wire_con_in_stage0[63]), .outData_64(wire_con_in_stage0[64]), .outData_65(wire_con_in_stage0[65]), .outData_66(wire_con_in_stage0[66]), .outData_67(wire_con_in_stage0[67]), .outData_68(wire_con_in_stage0[68]), .outData_69(wire_con_in_stage0[69]), .outData_70(wire_con_in_stage0[70]), .outData_71(wire_con_in_stage0[71]), .outData_72(wire_con_in_stage0[72]), .outData_73(wire_con_in_stage0[73]), .outData_74(wire_con_in_stage0[74]), .outData_75(wire_con_in_stage0[75]), .outData_76(wire_con_in_stage0[76]), .outData_77(wire_con_in_stage0[77]), .outData_78(wire_con_in_stage0[78]), .outData_79(wire_con_in_stage0[79]), .outData_80(wire_con_in_stage0[80]), .outData_81(wire_con_in_stage0[81]), .outData_82(wire_con_in_stage0[82]), .outData_83(wire_con_in_stage0[83]), .outData_84(wire_con_in_stage0[84]), .outData_85(wire_con_in_stage0[85]), .outData_86(wire_con_in_stage0[86]), .outData_87(wire_con_in_stage0[87]), .outData_88(wire_con_in_stage0[88]), .outData_89(wire_con_in_stage0[89]), .outData_90(wire_con_in_stage0[90]), .outData_91(wire_con_in_stage0[91]), .outData_92(wire_con_in_stage0[92]), .outData_93(wire_con_in_stage0[93]), .outData_94(wire_con_in_stage0[94]), .outData_95(wire_con_in_stage0[95]), .outData_96(wire_con_in_stage0[96]), .outData_97(wire_con_in_stage0[97]), .outData_98(wire_con_in_stage0[98]), .outData_99(wire_con_in_stage0[99]), .outData_100(wire_con_in_stage0[100]), .outData_101(wire_con_in_stage0[101]), .outData_102(wire_con_in_stage0[102]), .outData_103(wire_con_in_stage0[103]), .outData_104(wire_con_in_stage0[104]), .outData_105(wire_con_in_stage0[105]), .outData_106(wire_con_in_stage0[106]), .outData_107(wire_con_in_stage0[107]), .outData_108(wire_con_in_stage0[108]), .outData_109(wire_con_in_stage0[109]), .outData_110(wire_con_in_stage0[110]), .outData_111(wire_con_in_stage0[111]), .outData_112(wire_con_in_stage0[112]), .outData_113(wire_con_in_stage0[113]), .outData_114(wire_con_in_stage0[114]), .outData_115(wire_con_in_stage0[115]), .outData_116(wire_con_in_stage0[116]), .outData_117(wire_con_in_stage0[117]), .outData_118(wire_con_in_stage0[118]), .outData_119(wire_con_in_stage0[119]), .outData_120(wire_con_in_stage0[120]), .outData_121(wire_con_in_stage0[121]), .outData_122(wire_con_in_stage0[122]), .outData_123(wire_con_in_stage0[123]), .outData_124(wire_con_in_stage0[124]), .outData_125(wire_con_in_stage0[125]), .outData_126(wire_con_in_stage0[126]), .outData_127(wire_con_in_stage0[127]), .outData_128(wire_con_in_stage0[128]), .outData_129(wire_con_in_stage0[129]), .outData_130(wire_con_in_stage0[130]), .outData_131(wire_con_in_stage0[131]), .outData_132(wire_con_in_stage0[132]), .outData_133(wire_con_in_stage0[133]), .outData_134(wire_con_in_stage0[134]), .outData_135(wire_con_in_stage0[135]), .outData_136(wire_con_in_stage0[136]), .outData_137(wire_con_in_stage0[137]), .outData_138(wire_con_in_stage0[138]), .outData_139(wire_con_in_stage0[139]), .outData_140(wire_con_in_stage0[140]), .outData_141(wire_con_in_stage0[141]), .outData_142(wire_con_in_stage0[142]), .outData_143(wire_con_in_stage0[143]), .outData_144(wire_con_in_stage0[144]), .outData_145(wire_con_in_stage0[145]), .outData_146(wire_con_in_stage0[146]), .outData_147(wire_con_in_stage0[147]), .outData_148(wire_con_in_stage0[148]), .outData_149(wire_con_in_stage0[149]), .outData_150(wire_con_in_stage0[150]), .outData_151(wire_con_in_stage0[151]), .outData_152(wire_con_in_stage0[152]), .outData_153(wire_con_in_stage0[153]), .outData_154(wire_con_in_stage0[154]), .outData_155(wire_con_in_stage0[155]), .outData_156(wire_con_in_stage0[156]), .outData_157(wire_con_in_stage0[157]), .outData_158(wire_con_in_stage0[158]), .outData_159(wire_con_in_stage0[159]), .outData_160(wire_con_in_stage0[160]), .outData_161(wire_con_in_stage0[161]), .outData_162(wire_con_in_stage0[162]), .outData_163(wire_con_in_stage0[163]), .outData_164(wire_con_in_stage0[164]), .outData_165(wire_con_in_stage0[165]), .outData_166(wire_con_in_stage0[166]), .outData_167(wire_con_in_stage0[167]), .outData_168(wire_con_in_stage0[168]), .outData_169(wire_con_in_stage0[169]), .outData_170(wire_con_in_stage0[170]), .outData_171(wire_con_in_stage0[171]), .outData_172(wire_con_in_stage0[172]), .outData_173(wire_con_in_stage0[173]), .outData_174(wire_con_in_stage0[174]), .outData_175(wire_con_in_stage0[175]), .outData_176(wire_con_in_stage0[176]), .outData_177(wire_con_in_stage0[177]), .outData_178(wire_con_in_stage0[178]), .outData_179(wire_con_in_stage0[179]), .outData_180(wire_con_in_stage0[180]), .outData_181(wire_con_in_stage0[181]), .outData_182(wire_con_in_stage0[182]), .outData_183(wire_con_in_stage0[183]), .outData_184(wire_con_in_stage0[184]), .outData_185(wire_con_in_stage0[185]), .outData_186(wire_con_in_stage0[186]), .outData_187(wire_con_in_stage0[187]), .outData_188(wire_con_in_stage0[188]), .outData_189(wire_con_in_stage0[189]), .outData_190(wire_con_in_stage0[190]), .outData_191(wire_con_in_stage0[191]), .outData_192(wire_con_in_stage0[192]), .outData_193(wire_con_in_stage0[193]), .outData_194(wire_con_in_stage0[194]), .outData_195(wire_con_in_stage0[195]), .outData_196(wire_con_in_stage0[196]), .outData_197(wire_con_in_stage0[197]), .outData_198(wire_con_in_stage0[198]), .outData_199(wire_con_in_stage0[199]), .outData_200(wire_con_in_stage0[200]), .outData_201(wire_con_in_stage0[201]), .outData_202(wire_con_in_stage0[202]), .outData_203(wire_con_in_stage0[203]), .outData_204(wire_con_in_stage0[204]), .outData_205(wire_con_in_stage0[205]), .outData_206(wire_con_in_stage0[206]), .outData_207(wire_con_in_stage0[207]), .outData_208(wire_con_in_stage0[208]), .outData_209(wire_con_in_stage0[209]), .outData_210(wire_con_in_stage0[210]), .outData_211(wire_con_in_stage0[211]), .outData_212(wire_con_in_stage0[212]), .outData_213(wire_con_in_stage0[213]), .outData_214(wire_con_in_stage0[214]), .outData_215(wire_con_in_stage0[215]), .outData_216(wire_con_in_stage0[216]), .outData_217(wire_con_in_stage0[217]), .outData_218(wire_con_in_stage0[218]), .outData_219(wire_con_in_stage0[219]), .outData_220(wire_con_in_stage0[220]), .outData_221(wire_con_in_stage0[221]), .outData_222(wire_con_in_stage0[222]), .outData_223(wire_con_in_stage0[223]), .outData_224(wire_con_in_stage0[224]), .outData_225(wire_con_in_stage0[225]), .outData_226(wire_con_in_stage0[226]), .outData_227(wire_con_in_stage0[227]), .outData_228(wire_con_in_stage0[228]), .outData_229(wire_con_in_stage0[229]), .outData_230(wire_con_in_stage0[230]), .outData_231(wire_con_in_stage0[231]), .outData_232(wire_con_in_stage0[232]), .outData_233(wire_con_in_stage0[233]), .outData_234(wire_con_in_stage0[234]), .outData_235(wire_con_in_stage0[235]), .outData_236(wire_con_in_stage0[236]), .outData_237(wire_con_in_stage0[237]), .outData_238(wire_con_in_stage0[238]), .outData_239(wire_con_in_stage0[239]), .outData_240(wire_con_in_stage0[240]), .outData_241(wire_con_in_stage0[241]), .outData_242(wire_con_in_stage0[242]), .outData_243(wire_con_in_stage0[243]), .outData_244(wire_con_in_stage0[244]), .outData_245(wire_con_in_stage0[245]), .outData_246(wire_con_in_stage0[246]), .outData_247(wire_con_in_stage0[247]), .outData_248(wire_con_in_stage0[248]), .outData_249(wire_con_in_stage0[249]), .outData_250(wire_con_in_stage0[250]), .outData_251(wire_con_in_stage0[251]), .outData_252(wire_con_in_stage0[252]), .outData_253(wire_con_in_stage0[253]), .outData_254(wire_con_in_stage0[254]), .outData_255(wire_con_in_stage0[255]), 
        .in_start(in_start_stage0), .out_start(con_in_start_stage0), .ctrl(wire_ctrl_stage0), .clk(clk), .rst(rst));
  
  wireCon_dp256_st0_L wire_stage_0(
        .inData_0(wire_con_in_stage0[0]), .inData_1(wire_con_in_stage0[1]), .inData_2(wire_con_in_stage0[2]), .inData_3(wire_con_in_stage0[3]), .inData_4(wire_con_in_stage0[4]), .inData_5(wire_con_in_stage0[5]), .inData_6(wire_con_in_stage0[6]), .inData_7(wire_con_in_stage0[7]), .inData_8(wire_con_in_stage0[8]), .inData_9(wire_con_in_stage0[9]), .inData_10(wire_con_in_stage0[10]), .inData_11(wire_con_in_stage0[11]), .inData_12(wire_con_in_stage0[12]), .inData_13(wire_con_in_stage0[13]), .inData_14(wire_con_in_stage0[14]), .inData_15(wire_con_in_stage0[15]), .inData_16(wire_con_in_stage0[16]), .inData_17(wire_con_in_stage0[17]), .inData_18(wire_con_in_stage0[18]), .inData_19(wire_con_in_stage0[19]), .inData_20(wire_con_in_stage0[20]), .inData_21(wire_con_in_stage0[21]), .inData_22(wire_con_in_stage0[22]), .inData_23(wire_con_in_stage0[23]), .inData_24(wire_con_in_stage0[24]), .inData_25(wire_con_in_stage0[25]), .inData_26(wire_con_in_stage0[26]), .inData_27(wire_con_in_stage0[27]), .inData_28(wire_con_in_stage0[28]), .inData_29(wire_con_in_stage0[29]), .inData_30(wire_con_in_stage0[30]), .inData_31(wire_con_in_stage0[31]), .inData_32(wire_con_in_stage0[32]), .inData_33(wire_con_in_stage0[33]), .inData_34(wire_con_in_stage0[34]), .inData_35(wire_con_in_stage0[35]), .inData_36(wire_con_in_stage0[36]), .inData_37(wire_con_in_stage0[37]), .inData_38(wire_con_in_stage0[38]), .inData_39(wire_con_in_stage0[39]), .inData_40(wire_con_in_stage0[40]), .inData_41(wire_con_in_stage0[41]), .inData_42(wire_con_in_stage0[42]), .inData_43(wire_con_in_stage0[43]), .inData_44(wire_con_in_stage0[44]), .inData_45(wire_con_in_stage0[45]), .inData_46(wire_con_in_stage0[46]), .inData_47(wire_con_in_stage0[47]), .inData_48(wire_con_in_stage0[48]), .inData_49(wire_con_in_stage0[49]), .inData_50(wire_con_in_stage0[50]), .inData_51(wire_con_in_stage0[51]), .inData_52(wire_con_in_stage0[52]), .inData_53(wire_con_in_stage0[53]), .inData_54(wire_con_in_stage0[54]), .inData_55(wire_con_in_stage0[55]), .inData_56(wire_con_in_stage0[56]), .inData_57(wire_con_in_stage0[57]), .inData_58(wire_con_in_stage0[58]), .inData_59(wire_con_in_stage0[59]), .inData_60(wire_con_in_stage0[60]), .inData_61(wire_con_in_stage0[61]), .inData_62(wire_con_in_stage0[62]), .inData_63(wire_con_in_stage0[63]), .inData_64(wire_con_in_stage0[64]), .inData_65(wire_con_in_stage0[65]), .inData_66(wire_con_in_stage0[66]), .inData_67(wire_con_in_stage0[67]), .inData_68(wire_con_in_stage0[68]), .inData_69(wire_con_in_stage0[69]), .inData_70(wire_con_in_stage0[70]), .inData_71(wire_con_in_stage0[71]), .inData_72(wire_con_in_stage0[72]), .inData_73(wire_con_in_stage0[73]), .inData_74(wire_con_in_stage0[74]), .inData_75(wire_con_in_stage0[75]), .inData_76(wire_con_in_stage0[76]), .inData_77(wire_con_in_stage0[77]), .inData_78(wire_con_in_stage0[78]), .inData_79(wire_con_in_stage0[79]), .inData_80(wire_con_in_stage0[80]), .inData_81(wire_con_in_stage0[81]), .inData_82(wire_con_in_stage0[82]), .inData_83(wire_con_in_stage0[83]), .inData_84(wire_con_in_stage0[84]), .inData_85(wire_con_in_stage0[85]), .inData_86(wire_con_in_stage0[86]), .inData_87(wire_con_in_stage0[87]), .inData_88(wire_con_in_stage0[88]), .inData_89(wire_con_in_stage0[89]), .inData_90(wire_con_in_stage0[90]), .inData_91(wire_con_in_stage0[91]), .inData_92(wire_con_in_stage0[92]), .inData_93(wire_con_in_stage0[93]), .inData_94(wire_con_in_stage0[94]), .inData_95(wire_con_in_stage0[95]), .inData_96(wire_con_in_stage0[96]), .inData_97(wire_con_in_stage0[97]), .inData_98(wire_con_in_stage0[98]), .inData_99(wire_con_in_stage0[99]), .inData_100(wire_con_in_stage0[100]), .inData_101(wire_con_in_stage0[101]), .inData_102(wire_con_in_stage0[102]), .inData_103(wire_con_in_stage0[103]), .inData_104(wire_con_in_stage0[104]), .inData_105(wire_con_in_stage0[105]), .inData_106(wire_con_in_stage0[106]), .inData_107(wire_con_in_stage0[107]), .inData_108(wire_con_in_stage0[108]), .inData_109(wire_con_in_stage0[109]), .inData_110(wire_con_in_stage0[110]), .inData_111(wire_con_in_stage0[111]), .inData_112(wire_con_in_stage0[112]), .inData_113(wire_con_in_stage0[113]), .inData_114(wire_con_in_stage0[114]), .inData_115(wire_con_in_stage0[115]), .inData_116(wire_con_in_stage0[116]), .inData_117(wire_con_in_stage0[117]), .inData_118(wire_con_in_stage0[118]), .inData_119(wire_con_in_stage0[119]), .inData_120(wire_con_in_stage0[120]), .inData_121(wire_con_in_stage0[121]), .inData_122(wire_con_in_stage0[122]), .inData_123(wire_con_in_stage0[123]), .inData_124(wire_con_in_stage0[124]), .inData_125(wire_con_in_stage0[125]), .inData_126(wire_con_in_stage0[126]), .inData_127(wire_con_in_stage0[127]), .inData_128(wire_con_in_stage0[128]), .inData_129(wire_con_in_stage0[129]), .inData_130(wire_con_in_stage0[130]), .inData_131(wire_con_in_stage0[131]), .inData_132(wire_con_in_stage0[132]), .inData_133(wire_con_in_stage0[133]), .inData_134(wire_con_in_stage0[134]), .inData_135(wire_con_in_stage0[135]), .inData_136(wire_con_in_stage0[136]), .inData_137(wire_con_in_stage0[137]), .inData_138(wire_con_in_stage0[138]), .inData_139(wire_con_in_stage0[139]), .inData_140(wire_con_in_stage0[140]), .inData_141(wire_con_in_stage0[141]), .inData_142(wire_con_in_stage0[142]), .inData_143(wire_con_in_stage0[143]), .inData_144(wire_con_in_stage0[144]), .inData_145(wire_con_in_stage0[145]), .inData_146(wire_con_in_stage0[146]), .inData_147(wire_con_in_stage0[147]), .inData_148(wire_con_in_stage0[148]), .inData_149(wire_con_in_stage0[149]), .inData_150(wire_con_in_stage0[150]), .inData_151(wire_con_in_stage0[151]), .inData_152(wire_con_in_stage0[152]), .inData_153(wire_con_in_stage0[153]), .inData_154(wire_con_in_stage0[154]), .inData_155(wire_con_in_stage0[155]), .inData_156(wire_con_in_stage0[156]), .inData_157(wire_con_in_stage0[157]), .inData_158(wire_con_in_stage0[158]), .inData_159(wire_con_in_stage0[159]), .inData_160(wire_con_in_stage0[160]), .inData_161(wire_con_in_stage0[161]), .inData_162(wire_con_in_stage0[162]), .inData_163(wire_con_in_stage0[163]), .inData_164(wire_con_in_stage0[164]), .inData_165(wire_con_in_stage0[165]), .inData_166(wire_con_in_stage0[166]), .inData_167(wire_con_in_stage0[167]), .inData_168(wire_con_in_stage0[168]), .inData_169(wire_con_in_stage0[169]), .inData_170(wire_con_in_stage0[170]), .inData_171(wire_con_in_stage0[171]), .inData_172(wire_con_in_stage0[172]), .inData_173(wire_con_in_stage0[173]), .inData_174(wire_con_in_stage0[174]), .inData_175(wire_con_in_stage0[175]), .inData_176(wire_con_in_stage0[176]), .inData_177(wire_con_in_stage0[177]), .inData_178(wire_con_in_stage0[178]), .inData_179(wire_con_in_stage0[179]), .inData_180(wire_con_in_stage0[180]), .inData_181(wire_con_in_stage0[181]), .inData_182(wire_con_in_stage0[182]), .inData_183(wire_con_in_stage0[183]), .inData_184(wire_con_in_stage0[184]), .inData_185(wire_con_in_stage0[185]), .inData_186(wire_con_in_stage0[186]), .inData_187(wire_con_in_stage0[187]), .inData_188(wire_con_in_stage0[188]), .inData_189(wire_con_in_stage0[189]), .inData_190(wire_con_in_stage0[190]), .inData_191(wire_con_in_stage0[191]), .inData_192(wire_con_in_stage0[192]), .inData_193(wire_con_in_stage0[193]), .inData_194(wire_con_in_stage0[194]), .inData_195(wire_con_in_stage0[195]), .inData_196(wire_con_in_stage0[196]), .inData_197(wire_con_in_stage0[197]), .inData_198(wire_con_in_stage0[198]), .inData_199(wire_con_in_stage0[199]), .inData_200(wire_con_in_stage0[200]), .inData_201(wire_con_in_stage0[201]), .inData_202(wire_con_in_stage0[202]), .inData_203(wire_con_in_stage0[203]), .inData_204(wire_con_in_stage0[204]), .inData_205(wire_con_in_stage0[205]), .inData_206(wire_con_in_stage0[206]), .inData_207(wire_con_in_stage0[207]), .inData_208(wire_con_in_stage0[208]), .inData_209(wire_con_in_stage0[209]), .inData_210(wire_con_in_stage0[210]), .inData_211(wire_con_in_stage0[211]), .inData_212(wire_con_in_stage0[212]), .inData_213(wire_con_in_stage0[213]), .inData_214(wire_con_in_stage0[214]), .inData_215(wire_con_in_stage0[215]), .inData_216(wire_con_in_stage0[216]), .inData_217(wire_con_in_stage0[217]), .inData_218(wire_con_in_stage0[218]), .inData_219(wire_con_in_stage0[219]), .inData_220(wire_con_in_stage0[220]), .inData_221(wire_con_in_stage0[221]), .inData_222(wire_con_in_stage0[222]), .inData_223(wire_con_in_stage0[223]), .inData_224(wire_con_in_stage0[224]), .inData_225(wire_con_in_stage0[225]), .inData_226(wire_con_in_stage0[226]), .inData_227(wire_con_in_stage0[227]), .inData_228(wire_con_in_stage0[228]), .inData_229(wire_con_in_stage0[229]), .inData_230(wire_con_in_stage0[230]), .inData_231(wire_con_in_stage0[231]), .inData_232(wire_con_in_stage0[232]), .inData_233(wire_con_in_stage0[233]), .inData_234(wire_con_in_stage0[234]), .inData_235(wire_con_in_stage0[235]), .inData_236(wire_con_in_stage0[236]), .inData_237(wire_con_in_stage0[237]), .inData_238(wire_con_in_stage0[238]), .inData_239(wire_con_in_stage0[239]), .inData_240(wire_con_in_stage0[240]), .inData_241(wire_con_in_stage0[241]), .inData_242(wire_con_in_stage0[242]), .inData_243(wire_con_in_stage0[243]), .inData_244(wire_con_in_stage0[244]), .inData_245(wire_con_in_stage0[245]), .inData_246(wire_con_in_stage0[246]), .inData_247(wire_con_in_stage0[247]), .inData_248(wire_con_in_stage0[248]), .inData_249(wire_con_in_stage0[249]), .inData_250(wire_con_in_stage0[250]), .inData_251(wire_con_in_stage0[251]), .inData_252(wire_con_in_stage0[252]), .inData_253(wire_con_in_stage0[253]), .inData_254(wire_con_in_stage0[254]), .inData_255(wire_con_in_stage0[255]), 
        .outData_0(wire_con_out_stage0[0]), .outData_1(wire_con_out_stage0[1]), .outData_2(wire_con_out_stage0[2]), .outData_3(wire_con_out_stage0[3]), .outData_4(wire_con_out_stage0[4]), .outData_5(wire_con_out_stage0[5]), .outData_6(wire_con_out_stage0[6]), .outData_7(wire_con_out_stage0[7]), .outData_8(wire_con_out_stage0[8]), .outData_9(wire_con_out_stage0[9]), .outData_10(wire_con_out_stage0[10]), .outData_11(wire_con_out_stage0[11]), .outData_12(wire_con_out_stage0[12]), .outData_13(wire_con_out_stage0[13]), .outData_14(wire_con_out_stage0[14]), .outData_15(wire_con_out_stage0[15]), .outData_16(wire_con_out_stage0[16]), .outData_17(wire_con_out_stage0[17]), .outData_18(wire_con_out_stage0[18]), .outData_19(wire_con_out_stage0[19]), .outData_20(wire_con_out_stage0[20]), .outData_21(wire_con_out_stage0[21]), .outData_22(wire_con_out_stage0[22]), .outData_23(wire_con_out_stage0[23]), .outData_24(wire_con_out_stage0[24]), .outData_25(wire_con_out_stage0[25]), .outData_26(wire_con_out_stage0[26]), .outData_27(wire_con_out_stage0[27]), .outData_28(wire_con_out_stage0[28]), .outData_29(wire_con_out_stage0[29]), .outData_30(wire_con_out_stage0[30]), .outData_31(wire_con_out_stage0[31]), .outData_32(wire_con_out_stage0[32]), .outData_33(wire_con_out_stage0[33]), .outData_34(wire_con_out_stage0[34]), .outData_35(wire_con_out_stage0[35]), .outData_36(wire_con_out_stage0[36]), .outData_37(wire_con_out_stage0[37]), .outData_38(wire_con_out_stage0[38]), .outData_39(wire_con_out_stage0[39]), .outData_40(wire_con_out_stage0[40]), .outData_41(wire_con_out_stage0[41]), .outData_42(wire_con_out_stage0[42]), .outData_43(wire_con_out_stage0[43]), .outData_44(wire_con_out_stage0[44]), .outData_45(wire_con_out_stage0[45]), .outData_46(wire_con_out_stage0[46]), .outData_47(wire_con_out_stage0[47]), .outData_48(wire_con_out_stage0[48]), .outData_49(wire_con_out_stage0[49]), .outData_50(wire_con_out_stage0[50]), .outData_51(wire_con_out_stage0[51]), .outData_52(wire_con_out_stage0[52]), .outData_53(wire_con_out_stage0[53]), .outData_54(wire_con_out_stage0[54]), .outData_55(wire_con_out_stage0[55]), .outData_56(wire_con_out_stage0[56]), .outData_57(wire_con_out_stage0[57]), .outData_58(wire_con_out_stage0[58]), .outData_59(wire_con_out_stage0[59]), .outData_60(wire_con_out_stage0[60]), .outData_61(wire_con_out_stage0[61]), .outData_62(wire_con_out_stage0[62]), .outData_63(wire_con_out_stage0[63]), .outData_64(wire_con_out_stage0[64]), .outData_65(wire_con_out_stage0[65]), .outData_66(wire_con_out_stage0[66]), .outData_67(wire_con_out_stage0[67]), .outData_68(wire_con_out_stage0[68]), .outData_69(wire_con_out_stage0[69]), .outData_70(wire_con_out_stage0[70]), .outData_71(wire_con_out_stage0[71]), .outData_72(wire_con_out_stage0[72]), .outData_73(wire_con_out_stage0[73]), .outData_74(wire_con_out_stage0[74]), .outData_75(wire_con_out_stage0[75]), .outData_76(wire_con_out_stage0[76]), .outData_77(wire_con_out_stage0[77]), .outData_78(wire_con_out_stage0[78]), .outData_79(wire_con_out_stage0[79]), .outData_80(wire_con_out_stage0[80]), .outData_81(wire_con_out_stage0[81]), .outData_82(wire_con_out_stage0[82]), .outData_83(wire_con_out_stage0[83]), .outData_84(wire_con_out_stage0[84]), .outData_85(wire_con_out_stage0[85]), .outData_86(wire_con_out_stage0[86]), .outData_87(wire_con_out_stage0[87]), .outData_88(wire_con_out_stage0[88]), .outData_89(wire_con_out_stage0[89]), .outData_90(wire_con_out_stage0[90]), .outData_91(wire_con_out_stage0[91]), .outData_92(wire_con_out_stage0[92]), .outData_93(wire_con_out_stage0[93]), .outData_94(wire_con_out_stage0[94]), .outData_95(wire_con_out_stage0[95]), .outData_96(wire_con_out_stage0[96]), .outData_97(wire_con_out_stage0[97]), .outData_98(wire_con_out_stage0[98]), .outData_99(wire_con_out_stage0[99]), .outData_100(wire_con_out_stage0[100]), .outData_101(wire_con_out_stage0[101]), .outData_102(wire_con_out_stage0[102]), .outData_103(wire_con_out_stage0[103]), .outData_104(wire_con_out_stage0[104]), .outData_105(wire_con_out_stage0[105]), .outData_106(wire_con_out_stage0[106]), .outData_107(wire_con_out_stage0[107]), .outData_108(wire_con_out_stage0[108]), .outData_109(wire_con_out_stage0[109]), .outData_110(wire_con_out_stage0[110]), .outData_111(wire_con_out_stage0[111]), .outData_112(wire_con_out_stage0[112]), .outData_113(wire_con_out_stage0[113]), .outData_114(wire_con_out_stage0[114]), .outData_115(wire_con_out_stage0[115]), .outData_116(wire_con_out_stage0[116]), .outData_117(wire_con_out_stage0[117]), .outData_118(wire_con_out_stage0[118]), .outData_119(wire_con_out_stage0[119]), .outData_120(wire_con_out_stage0[120]), .outData_121(wire_con_out_stage0[121]), .outData_122(wire_con_out_stage0[122]), .outData_123(wire_con_out_stage0[123]), .outData_124(wire_con_out_stage0[124]), .outData_125(wire_con_out_stage0[125]), .outData_126(wire_con_out_stage0[126]), .outData_127(wire_con_out_stage0[127]), .outData_128(wire_con_out_stage0[128]), .outData_129(wire_con_out_stage0[129]), .outData_130(wire_con_out_stage0[130]), .outData_131(wire_con_out_stage0[131]), .outData_132(wire_con_out_stage0[132]), .outData_133(wire_con_out_stage0[133]), .outData_134(wire_con_out_stage0[134]), .outData_135(wire_con_out_stage0[135]), .outData_136(wire_con_out_stage0[136]), .outData_137(wire_con_out_stage0[137]), .outData_138(wire_con_out_stage0[138]), .outData_139(wire_con_out_stage0[139]), .outData_140(wire_con_out_stage0[140]), .outData_141(wire_con_out_stage0[141]), .outData_142(wire_con_out_stage0[142]), .outData_143(wire_con_out_stage0[143]), .outData_144(wire_con_out_stage0[144]), .outData_145(wire_con_out_stage0[145]), .outData_146(wire_con_out_stage0[146]), .outData_147(wire_con_out_stage0[147]), .outData_148(wire_con_out_stage0[148]), .outData_149(wire_con_out_stage0[149]), .outData_150(wire_con_out_stage0[150]), .outData_151(wire_con_out_stage0[151]), .outData_152(wire_con_out_stage0[152]), .outData_153(wire_con_out_stage0[153]), .outData_154(wire_con_out_stage0[154]), .outData_155(wire_con_out_stage0[155]), .outData_156(wire_con_out_stage0[156]), .outData_157(wire_con_out_stage0[157]), .outData_158(wire_con_out_stage0[158]), .outData_159(wire_con_out_stage0[159]), .outData_160(wire_con_out_stage0[160]), .outData_161(wire_con_out_stage0[161]), .outData_162(wire_con_out_stage0[162]), .outData_163(wire_con_out_stage0[163]), .outData_164(wire_con_out_stage0[164]), .outData_165(wire_con_out_stage0[165]), .outData_166(wire_con_out_stage0[166]), .outData_167(wire_con_out_stage0[167]), .outData_168(wire_con_out_stage0[168]), .outData_169(wire_con_out_stage0[169]), .outData_170(wire_con_out_stage0[170]), .outData_171(wire_con_out_stage0[171]), .outData_172(wire_con_out_stage0[172]), .outData_173(wire_con_out_stage0[173]), .outData_174(wire_con_out_stage0[174]), .outData_175(wire_con_out_stage0[175]), .outData_176(wire_con_out_stage0[176]), .outData_177(wire_con_out_stage0[177]), .outData_178(wire_con_out_stage0[178]), .outData_179(wire_con_out_stage0[179]), .outData_180(wire_con_out_stage0[180]), .outData_181(wire_con_out_stage0[181]), .outData_182(wire_con_out_stage0[182]), .outData_183(wire_con_out_stage0[183]), .outData_184(wire_con_out_stage0[184]), .outData_185(wire_con_out_stage0[185]), .outData_186(wire_con_out_stage0[186]), .outData_187(wire_con_out_stage0[187]), .outData_188(wire_con_out_stage0[188]), .outData_189(wire_con_out_stage0[189]), .outData_190(wire_con_out_stage0[190]), .outData_191(wire_con_out_stage0[191]), .outData_192(wire_con_out_stage0[192]), .outData_193(wire_con_out_stage0[193]), .outData_194(wire_con_out_stage0[194]), .outData_195(wire_con_out_stage0[195]), .outData_196(wire_con_out_stage0[196]), .outData_197(wire_con_out_stage0[197]), .outData_198(wire_con_out_stage0[198]), .outData_199(wire_con_out_stage0[199]), .outData_200(wire_con_out_stage0[200]), .outData_201(wire_con_out_stage0[201]), .outData_202(wire_con_out_stage0[202]), .outData_203(wire_con_out_stage0[203]), .outData_204(wire_con_out_stage0[204]), .outData_205(wire_con_out_stage0[205]), .outData_206(wire_con_out_stage0[206]), .outData_207(wire_con_out_stage0[207]), .outData_208(wire_con_out_stage0[208]), .outData_209(wire_con_out_stage0[209]), .outData_210(wire_con_out_stage0[210]), .outData_211(wire_con_out_stage0[211]), .outData_212(wire_con_out_stage0[212]), .outData_213(wire_con_out_stage0[213]), .outData_214(wire_con_out_stage0[214]), .outData_215(wire_con_out_stage0[215]), .outData_216(wire_con_out_stage0[216]), .outData_217(wire_con_out_stage0[217]), .outData_218(wire_con_out_stage0[218]), .outData_219(wire_con_out_stage0[219]), .outData_220(wire_con_out_stage0[220]), .outData_221(wire_con_out_stage0[221]), .outData_222(wire_con_out_stage0[222]), .outData_223(wire_con_out_stage0[223]), .outData_224(wire_con_out_stage0[224]), .outData_225(wire_con_out_stage0[225]), .outData_226(wire_con_out_stage0[226]), .outData_227(wire_con_out_stage0[227]), .outData_228(wire_con_out_stage0[228]), .outData_229(wire_con_out_stage0[229]), .outData_230(wire_con_out_stage0[230]), .outData_231(wire_con_out_stage0[231]), .outData_232(wire_con_out_stage0[232]), .outData_233(wire_con_out_stage0[233]), .outData_234(wire_con_out_stage0[234]), .outData_235(wire_con_out_stage0[235]), .outData_236(wire_con_out_stage0[236]), .outData_237(wire_con_out_stage0[237]), .outData_238(wire_con_out_stage0[238]), .outData_239(wire_con_out_stage0[239]), .outData_240(wire_con_out_stage0[240]), .outData_241(wire_con_out_stage0[241]), .outData_242(wire_con_out_stage0[242]), .outData_243(wire_con_out_stage0[243]), .outData_244(wire_con_out_stage0[244]), .outData_245(wire_con_out_stage0[245]), .outData_246(wire_con_out_stage0[246]), .outData_247(wire_con_out_stage0[247]), .outData_248(wire_con_out_stage0[248]), .outData_249(wire_con_out_stage0[249]), .outData_250(wire_con_out_stage0[250]), .outData_251(wire_con_out_stage0[251]), .outData_252(wire_con_out_stage0[252]), .outData_253(wire_con_out_stage0[253]), .outData_254(wire_con_out_stage0[254]), .outData_255(wire_con_out_stage0[255]), 
        .in_start(con_in_start_stage0), .out_start(in_start_stage1), .clk(clk), .rst(rst)); 

  
  wire [7:0] counter_w;
  assign counter_w = counter_in; 
  assign wire_ctrl_stage0[0] = counter_w[7]; 
  assign wire_ctrl_stage0[1] = counter_w[7]; 
  assign wire_ctrl_stage0[2] = counter_w[7]; 
  assign wire_ctrl_stage0[3] = counter_w[7]; 
  assign wire_ctrl_stage0[4] = counter_w[7]; 
  assign wire_ctrl_stage0[5] = counter_w[7]; 
  assign wire_ctrl_stage0[6] = counter_w[7]; 
  assign wire_ctrl_stage0[7] = counter_w[7]; 
  assign wire_ctrl_stage0[8] = counter_w[7]; 
  assign wire_ctrl_stage0[9] = counter_w[7]; 
  assign wire_ctrl_stage0[10] = counter_w[7]; 
  assign wire_ctrl_stage0[11] = counter_w[7]; 
  assign wire_ctrl_stage0[12] = counter_w[7]; 
  assign wire_ctrl_stage0[13] = counter_w[7]; 
  assign wire_ctrl_stage0[14] = counter_w[7]; 
  assign wire_ctrl_stage0[15] = counter_w[7]; 
  assign wire_ctrl_stage0[16] = counter_w[7]; 
  assign wire_ctrl_stage0[17] = counter_w[7]; 
  assign wire_ctrl_stage0[18] = counter_w[7]; 
  assign wire_ctrl_stage0[19] = counter_w[7]; 
  assign wire_ctrl_stage0[20] = counter_w[7]; 
  assign wire_ctrl_stage0[21] = counter_w[7]; 
  assign wire_ctrl_stage0[22] = counter_w[7]; 
  assign wire_ctrl_stage0[23] = counter_w[7]; 
  assign wire_ctrl_stage0[24] = counter_w[7]; 
  assign wire_ctrl_stage0[25] = counter_w[7]; 
  assign wire_ctrl_stage0[26] = counter_w[7]; 
  assign wire_ctrl_stage0[27] = counter_w[7]; 
  assign wire_ctrl_stage0[28] = counter_w[7]; 
  assign wire_ctrl_stage0[29] = counter_w[7]; 
  assign wire_ctrl_stage0[30] = counter_w[7]; 
  assign wire_ctrl_stage0[31] = counter_w[7]; 
  assign wire_ctrl_stage0[32] = counter_w[7]; 
  assign wire_ctrl_stage0[33] = counter_w[7]; 
  assign wire_ctrl_stage0[34] = counter_w[7]; 
  assign wire_ctrl_stage0[35] = counter_w[7]; 
  assign wire_ctrl_stage0[36] = counter_w[7]; 
  assign wire_ctrl_stage0[37] = counter_w[7]; 
  assign wire_ctrl_stage0[38] = counter_w[7]; 
  assign wire_ctrl_stage0[39] = counter_w[7]; 
  assign wire_ctrl_stage0[40] = counter_w[7]; 
  assign wire_ctrl_stage0[41] = counter_w[7]; 
  assign wire_ctrl_stage0[42] = counter_w[7]; 
  assign wire_ctrl_stage0[43] = counter_w[7]; 
  assign wire_ctrl_stage0[44] = counter_w[7]; 
  assign wire_ctrl_stage0[45] = counter_w[7]; 
  assign wire_ctrl_stage0[46] = counter_w[7]; 
  assign wire_ctrl_stage0[47] = counter_w[7]; 
  assign wire_ctrl_stage0[48] = counter_w[7]; 
  assign wire_ctrl_stage0[49] = counter_w[7]; 
  assign wire_ctrl_stage0[50] = counter_w[7]; 
  assign wire_ctrl_stage0[51] = counter_w[7]; 
  assign wire_ctrl_stage0[52] = counter_w[7]; 
  assign wire_ctrl_stage0[53] = counter_w[7]; 
  assign wire_ctrl_stage0[54] = counter_w[7]; 
  assign wire_ctrl_stage0[55] = counter_w[7]; 
  assign wire_ctrl_stage0[56] = counter_w[7]; 
  assign wire_ctrl_stage0[57] = counter_w[7]; 
  assign wire_ctrl_stage0[58] = counter_w[7]; 
  assign wire_ctrl_stage0[59] = counter_w[7]; 
  assign wire_ctrl_stage0[60] = counter_w[7]; 
  assign wire_ctrl_stage0[61] = counter_w[7]; 
  assign wire_ctrl_stage0[62] = counter_w[7]; 
  assign wire_ctrl_stage0[63] = counter_w[7]; 
  assign wire_ctrl_stage0[64] = counter_w[7]; 
  assign wire_ctrl_stage0[65] = counter_w[7]; 
  assign wire_ctrl_stage0[66] = counter_w[7]; 
  assign wire_ctrl_stage0[67] = counter_w[7]; 
  assign wire_ctrl_stage0[68] = counter_w[7]; 
  assign wire_ctrl_stage0[69] = counter_w[7]; 
  assign wire_ctrl_stage0[70] = counter_w[7]; 
  assign wire_ctrl_stage0[71] = counter_w[7]; 
  assign wire_ctrl_stage0[72] = counter_w[7]; 
  assign wire_ctrl_stage0[73] = counter_w[7]; 
  assign wire_ctrl_stage0[74] = counter_w[7]; 
  assign wire_ctrl_stage0[75] = counter_w[7]; 
  assign wire_ctrl_stage0[76] = counter_w[7]; 
  assign wire_ctrl_stage0[77] = counter_w[7]; 
  assign wire_ctrl_stage0[78] = counter_w[7]; 
  assign wire_ctrl_stage0[79] = counter_w[7]; 
  assign wire_ctrl_stage0[80] = counter_w[7]; 
  assign wire_ctrl_stage0[81] = counter_w[7]; 
  assign wire_ctrl_stage0[82] = counter_w[7]; 
  assign wire_ctrl_stage0[83] = counter_w[7]; 
  assign wire_ctrl_stage0[84] = counter_w[7]; 
  assign wire_ctrl_stage0[85] = counter_w[7]; 
  assign wire_ctrl_stage0[86] = counter_w[7]; 
  assign wire_ctrl_stage0[87] = counter_w[7]; 
  assign wire_ctrl_stage0[88] = counter_w[7]; 
  assign wire_ctrl_stage0[89] = counter_w[7]; 
  assign wire_ctrl_stage0[90] = counter_w[7]; 
  assign wire_ctrl_stage0[91] = counter_w[7]; 
  assign wire_ctrl_stage0[92] = counter_w[7]; 
  assign wire_ctrl_stage0[93] = counter_w[7]; 
  assign wire_ctrl_stage0[94] = counter_w[7]; 
  assign wire_ctrl_stage0[95] = counter_w[7]; 
  assign wire_ctrl_stage0[96] = counter_w[7]; 
  assign wire_ctrl_stage0[97] = counter_w[7]; 
  assign wire_ctrl_stage0[98] = counter_w[7]; 
  assign wire_ctrl_stage0[99] = counter_w[7]; 
  assign wire_ctrl_stage0[100] = counter_w[7]; 
  assign wire_ctrl_stage0[101] = counter_w[7]; 
  assign wire_ctrl_stage0[102] = counter_w[7]; 
  assign wire_ctrl_stage0[103] = counter_w[7]; 
  assign wire_ctrl_stage0[104] = counter_w[7]; 
  assign wire_ctrl_stage0[105] = counter_w[7]; 
  assign wire_ctrl_stage0[106] = counter_w[7]; 
  assign wire_ctrl_stage0[107] = counter_w[7]; 
  assign wire_ctrl_stage0[108] = counter_w[7]; 
  assign wire_ctrl_stage0[109] = counter_w[7]; 
  assign wire_ctrl_stage0[110] = counter_w[7]; 
  assign wire_ctrl_stage0[111] = counter_w[7]; 
  assign wire_ctrl_stage0[112] = counter_w[7]; 
  assign wire_ctrl_stage0[113] = counter_w[7]; 
  assign wire_ctrl_stage0[114] = counter_w[7]; 
  assign wire_ctrl_stage0[115] = counter_w[7]; 
  assign wire_ctrl_stage0[116] = counter_w[7]; 
  assign wire_ctrl_stage0[117] = counter_w[7]; 
  assign wire_ctrl_stage0[118] = counter_w[7]; 
  assign wire_ctrl_stage0[119] = counter_w[7]; 
  assign wire_ctrl_stage0[120] = counter_w[7]; 
  assign wire_ctrl_stage0[121] = counter_w[7]; 
  assign wire_ctrl_stage0[122] = counter_w[7]; 
  assign wire_ctrl_stage0[123] = counter_w[7]; 
  assign wire_ctrl_stage0[124] = counter_w[7]; 
  assign wire_ctrl_stage0[125] = counter_w[7]; 
  assign wire_ctrl_stage0[126] = counter_w[7]; 
  assign wire_ctrl_stage0[127] = counter_w[7]; 
  wire [DATA_WIDTH-1:0] wire_con_in_stage1[255:0];
  wire [DATA_WIDTH-1:0] wire_con_out_stage1[255:0];
  wire [127:0] wire_ctrl_stage1;

  switches_stage_st1_0_L switch_stage_1(
        .inData_0(wire_con_out_stage0[0]), .inData_1(wire_con_out_stage0[1]), .inData_2(wire_con_out_stage0[2]), .inData_3(wire_con_out_stage0[3]), .inData_4(wire_con_out_stage0[4]), .inData_5(wire_con_out_stage0[5]), .inData_6(wire_con_out_stage0[6]), .inData_7(wire_con_out_stage0[7]), .inData_8(wire_con_out_stage0[8]), .inData_9(wire_con_out_stage0[9]), .inData_10(wire_con_out_stage0[10]), .inData_11(wire_con_out_stage0[11]), .inData_12(wire_con_out_stage0[12]), .inData_13(wire_con_out_stage0[13]), .inData_14(wire_con_out_stage0[14]), .inData_15(wire_con_out_stage0[15]), .inData_16(wire_con_out_stage0[16]), .inData_17(wire_con_out_stage0[17]), .inData_18(wire_con_out_stage0[18]), .inData_19(wire_con_out_stage0[19]), .inData_20(wire_con_out_stage0[20]), .inData_21(wire_con_out_stage0[21]), .inData_22(wire_con_out_stage0[22]), .inData_23(wire_con_out_stage0[23]), .inData_24(wire_con_out_stage0[24]), .inData_25(wire_con_out_stage0[25]), .inData_26(wire_con_out_stage0[26]), .inData_27(wire_con_out_stage0[27]), .inData_28(wire_con_out_stage0[28]), .inData_29(wire_con_out_stage0[29]), .inData_30(wire_con_out_stage0[30]), .inData_31(wire_con_out_stage0[31]), .inData_32(wire_con_out_stage0[32]), .inData_33(wire_con_out_stage0[33]), .inData_34(wire_con_out_stage0[34]), .inData_35(wire_con_out_stage0[35]), .inData_36(wire_con_out_stage0[36]), .inData_37(wire_con_out_stage0[37]), .inData_38(wire_con_out_stage0[38]), .inData_39(wire_con_out_stage0[39]), .inData_40(wire_con_out_stage0[40]), .inData_41(wire_con_out_stage0[41]), .inData_42(wire_con_out_stage0[42]), .inData_43(wire_con_out_stage0[43]), .inData_44(wire_con_out_stage0[44]), .inData_45(wire_con_out_stage0[45]), .inData_46(wire_con_out_stage0[46]), .inData_47(wire_con_out_stage0[47]), .inData_48(wire_con_out_stage0[48]), .inData_49(wire_con_out_stage0[49]), .inData_50(wire_con_out_stage0[50]), .inData_51(wire_con_out_stage0[51]), .inData_52(wire_con_out_stage0[52]), .inData_53(wire_con_out_stage0[53]), .inData_54(wire_con_out_stage0[54]), .inData_55(wire_con_out_stage0[55]), .inData_56(wire_con_out_stage0[56]), .inData_57(wire_con_out_stage0[57]), .inData_58(wire_con_out_stage0[58]), .inData_59(wire_con_out_stage0[59]), .inData_60(wire_con_out_stage0[60]), .inData_61(wire_con_out_stage0[61]), .inData_62(wire_con_out_stage0[62]), .inData_63(wire_con_out_stage0[63]), .inData_64(wire_con_out_stage0[64]), .inData_65(wire_con_out_stage0[65]), .inData_66(wire_con_out_stage0[66]), .inData_67(wire_con_out_stage0[67]), .inData_68(wire_con_out_stage0[68]), .inData_69(wire_con_out_stage0[69]), .inData_70(wire_con_out_stage0[70]), .inData_71(wire_con_out_stage0[71]), .inData_72(wire_con_out_stage0[72]), .inData_73(wire_con_out_stage0[73]), .inData_74(wire_con_out_stage0[74]), .inData_75(wire_con_out_stage0[75]), .inData_76(wire_con_out_stage0[76]), .inData_77(wire_con_out_stage0[77]), .inData_78(wire_con_out_stage0[78]), .inData_79(wire_con_out_stage0[79]), .inData_80(wire_con_out_stage0[80]), .inData_81(wire_con_out_stage0[81]), .inData_82(wire_con_out_stage0[82]), .inData_83(wire_con_out_stage0[83]), .inData_84(wire_con_out_stage0[84]), .inData_85(wire_con_out_stage0[85]), .inData_86(wire_con_out_stage0[86]), .inData_87(wire_con_out_stage0[87]), .inData_88(wire_con_out_stage0[88]), .inData_89(wire_con_out_stage0[89]), .inData_90(wire_con_out_stage0[90]), .inData_91(wire_con_out_stage0[91]), .inData_92(wire_con_out_stage0[92]), .inData_93(wire_con_out_stage0[93]), .inData_94(wire_con_out_stage0[94]), .inData_95(wire_con_out_stage0[95]), .inData_96(wire_con_out_stage0[96]), .inData_97(wire_con_out_stage0[97]), .inData_98(wire_con_out_stage0[98]), .inData_99(wire_con_out_stage0[99]), .inData_100(wire_con_out_stage0[100]), .inData_101(wire_con_out_stage0[101]), .inData_102(wire_con_out_stage0[102]), .inData_103(wire_con_out_stage0[103]), .inData_104(wire_con_out_stage0[104]), .inData_105(wire_con_out_stage0[105]), .inData_106(wire_con_out_stage0[106]), .inData_107(wire_con_out_stage0[107]), .inData_108(wire_con_out_stage0[108]), .inData_109(wire_con_out_stage0[109]), .inData_110(wire_con_out_stage0[110]), .inData_111(wire_con_out_stage0[111]), .inData_112(wire_con_out_stage0[112]), .inData_113(wire_con_out_stage0[113]), .inData_114(wire_con_out_stage0[114]), .inData_115(wire_con_out_stage0[115]), .inData_116(wire_con_out_stage0[116]), .inData_117(wire_con_out_stage0[117]), .inData_118(wire_con_out_stage0[118]), .inData_119(wire_con_out_stage0[119]), .inData_120(wire_con_out_stage0[120]), .inData_121(wire_con_out_stage0[121]), .inData_122(wire_con_out_stage0[122]), .inData_123(wire_con_out_stage0[123]), .inData_124(wire_con_out_stage0[124]), .inData_125(wire_con_out_stage0[125]), .inData_126(wire_con_out_stage0[126]), .inData_127(wire_con_out_stage0[127]), .inData_128(wire_con_out_stage0[128]), .inData_129(wire_con_out_stage0[129]), .inData_130(wire_con_out_stage0[130]), .inData_131(wire_con_out_stage0[131]), .inData_132(wire_con_out_stage0[132]), .inData_133(wire_con_out_stage0[133]), .inData_134(wire_con_out_stage0[134]), .inData_135(wire_con_out_stage0[135]), .inData_136(wire_con_out_stage0[136]), .inData_137(wire_con_out_stage0[137]), .inData_138(wire_con_out_stage0[138]), .inData_139(wire_con_out_stage0[139]), .inData_140(wire_con_out_stage0[140]), .inData_141(wire_con_out_stage0[141]), .inData_142(wire_con_out_stage0[142]), .inData_143(wire_con_out_stage0[143]), .inData_144(wire_con_out_stage0[144]), .inData_145(wire_con_out_stage0[145]), .inData_146(wire_con_out_stage0[146]), .inData_147(wire_con_out_stage0[147]), .inData_148(wire_con_out_stage0[148]), .inData_149(wire_con_out_stage0[149]), .inData_150(wire_con_out_stage0[150]), .inData_151(wire_con_out_stage0[151]), .inData_152(wire_con_out_stage0[152]), .inData_153(wire_con_out_stage0[153]), .inData_154(wire_con_out_stage0[154]), .inData_155(wire_con_out_stage0[155]), .inData_156(wire_con_out_stage0[156]), .inData_157(wire_con_out_stage0[157]), .inData_158(wire_con_out_stage0[158]), .inData_159(wire_con_out_stage0[159]), .inData_160(wire_con_out_stage0[160]), .inData_161(wire_con_out_stage0[161]), .inData_162(wire_con_out_stage0[162]), .inData_163(wire_con_out_stage0[163]), .inData_164(wire_con_out_stage0[164]), .inData_165(wire_con_out_stage0[165]), .inData_166(wire_con_out_stage0[166]), .inData_167(wire_con_out_stage0[167]), .inData_168(wire_con_out_stage0[168]), .inData_169(wire_con_out_stage0[169]), .inData_170(wire_con_out_stage0[170]), .inData_171(wire_con_out_stage0[171]), .inData_172(wire_con_out_stage0[172]), .inData_173(wire_con_out_stage0[173]), .inData_174(wire_con_out_stage0[174]), .inData_175(wire_con_out_stage0[175]), .inData_176(wire_con_out_stage0[176]), .inData_177(wire_con_out_stage0[177]), .inData_178(wire_con_out_stage0[178]), .inData_179(wire_con_out_stage0[179]), .inData_180(wire_con_out_stage0[180]), .inData_181(wire_con_out_stage0[181]), .inData_182(wire_con_out_stage0[182]), .inData_183(wire_con_out_stage0[183]), .inData_184(wire_con_out_stage0[184]), .inData_185(wire_con_out_stage0[185]), .inData_186(wire_con_out_stage0[186]), .inData_187(wire_con_out_stage0[187]), .inData_188(wire_con_out_stage0[188]), .inData_189(wire_con_out_stage0[189]), .inData_190(wire_con_out_stage0[190]), .inData_191(wire_con_out_stage0[191]), .inData_192(wire_con_out_stage0[192]), .inData_193(wire_con_out_stage0[193]), .inData_194(wire_con_out_stage0[194]), .inData_195(wire_con_out_stage0[195]), .inData_196(wire_con_out_stage0[196]), .inData_197(wire_con_out_stage0[197]), .inData_198(wire_con_out_stage0[198]), .inData_199(wire_con_out_stage0[199]), .inData_200(wire_con_out_stage0[200]), .inData_201(wire_con_out_stage0[201]), .inData_202(wire_con_out_stage0[202]), .inData_203(wire_con_out_stage0[203]), .inData_204(wire_con_out_stage0[204]), .inData_205(wire_con_out_stage0[205]), .inData_206(wire_con_out_stage0[206]), .inData_207(wire_con_out_stage0[207]), .inData_208(wire_con_out_stage0[208]), .inData_209(wire_con_out_stage0[209]), .inData_210(wire_con_out_stage0[210]), .inData_211(wire_con_out_stage0[211]), .inData_212(wire_con_out_stage0[212]), .inData_213(wire_con_out_stage0[213]), .inData_214(wire_con_out_stage0[214]), .inData_215(wire_con_out_stage0[215]), .inData_216(wire_con_out_stage0[216]), .inData_217(wire_con_out_stage0[217]), .inData_218(wire_con_out_stage0[218]), .inData_219(wire_con_out_stage0[219]), .inData_220(wire_con_out_stage0[220]), .inData_221(wire_con_out_stage0[221]), .inData_222(wire_con_out_stage0[222]), .inData_223(wire_con_out_stage0[223]), .inData_224(wire_con_out_stage0[224]), .inData_225(wire_con_out_stage0[225]), .inData_226(wire_con_out_stage0[226]), .inData_227(wire_con_out_stage0[227]), .inData_228(wire_con_out_stage0[228]), .inData_229(wire_con_out_stage0[229]), .inData_230(wire_con_out_stage0[230]), .inData_231(wire_con_out_stage0[231]), .inData_232(wire_con_out_stage0[232]), .inData_233(wire_con_out_stage0[233]), .inData_234(wire_con_out_stage0[234]), .inData_235(wire_con_out_stage0[235]), .inData_236(wire_con_out_stage0[236]), .inData_237(wire_con_out_stage0[237]), .inData_238(wire_con_out_stage0[238]), .inData_239(wire_con_out_stage0[239]), .inData_240(wire_con_out_stage0[240]), .inData_241(wire_con_out_stage0[241]), .inData_242(wire_con_out_stage0[242]), .inData_243(wire_con_out_stage0[243]), .inData_244(wire_con_out_stage0[244]), .inData_245(wire_con_out_stage0[245]), .inData_246(wire_con_out_stage0[246]), .inData_247(wire_con_out_stage0[247]), .inData_248(wire_con_out_stage0[248]), .inData_249(wire_con_out_stage0[249]), .inData_250(wire_con_out_stage0[250]), .inData_251(wire_con_out_stage0[251]), .inData_252(wire_con_out_stage0[252]), .inData_253(wire_con_out_stage0[253]), .inData_254(wire_con_out_stage0[254]), .inData_255(wire_con_out_stage0[255]), 
        .outData_0(wire_con_in_stage1[0]), .outData_1(wire_con_in_stage1[1]), .outData_2(wire_con_in_stage1[2]), .outData_3(wire_con_in_stage1[3]), .outData_4(wire_con_in_stage1[4]), .outData_5(wire_con_in_stage1[5]), .outData_6(wire_con_in_stage1[6]), .outData_7(wire_con_in_stage1[7]), .outData_8(wire_con_in_stage1[8]), .outData_9(wire_con_in_stage1[9]), .outData_10(wire_con_in_stage1[10]), .outData_11(wire_con_in_stage1[11]), .outData_12(wire_con_in_stage1[12]), .outData_13(wire_con_in_stage1[13]), .outData_14(wire_con_in_stage1[14]), .outData_15(wire_con_in_stage1[15]), .outData_16(wire_con_in_stage1[16]), .outData_17(wire_con_in_stage1[17]), .outData_18(wire_con_in_stage1[18]), .outData_19(wire_con_in_stage1[19]), .outData_20(wire_con_in_stage1[20]), .outData_21(wire_con_in_stage1[21]), .outData_22(wire_con_in_stage1[22]), .outData_23(wire_con_in_stage1[23]), .outData_24(wire_con_in_stage1[24]), .outData_25(wire_con_in_stage1[25]), .outData_26(wire_con_in_stage1[26]), .outData_27(wire_con_in_stage1[27]), .outData_28(wire_con_in_stage1[28]), .outData_29(wire_con_in_stage1[29]), .outData_30(wire_con_in_stage1[30]), .outData_31(wire_con_in_stage1[31]), .outData_32(wire_con_in_stage1[32]), .outData_33(wire_con_in_stage1[33]), .outData_34(wire_con_in_stage1[34]), .outData_35(wire_con_in_stage1[35]), .outData_36(wire_con_in_stage1[36]), .outData_37(wire_con_in_stage1[37]), .outData_38(wire_con_in_stage1[38]), .outData_39(wire_con_in_stage1[39]), .outData_40(wire_con_in_stage1[40]), .outData_41(wire_con_in_stage1[41]), .outData_42(wire_con_in_stage1[42]), .outData_43(wire_con_in_stage1[43]), .outData_44(wire_con_in_stage1[44]), .outData_45(wire_con_in_stage1[45]), .outData_46(wire_con_in_stage1[46]), .outData_47(wire_con_in_stage1[47]), .outData_48(wire_con_in_stage1[48]), .outData_49(wire_con_in_stage1[49]), .outData_50(wire_con_in_stage1[50]), .outData_51(wire_con_in_stage1[51]), .outData_52(wire_con_in_stage1[52]), .outData_53(wire_con_in_stage1[53]), .outData_54(wire_con_in_stage1[54]), .outData_55(wire_con_in_stage1[55]), .outData_56(wire_con_in_stage1[56]), .outData_57(wire_con_in_stage1[57]), .outData_58(wire_con_in_stage1[58]), .outData_59(wire_con_in_stage1[59]), .outData_60(wire_con_in_stage1[60]), .outData_61(wire_con_in_stage1[61]), .outData_62(wire_con_in_stage1[62]), .outData_63(wire_con_in_stage1[63]), .outData_64(wire_con_in_stage1[64]), .outData_65(wire_con_in_stage1[65]), .outData_66(wire_con_in_stage1[66]), .outData_67(wire_con_in_stage1[67]), .outData_68(wire_con_in_stage1[68]), .outData_69(wire_con_in_stage1[69]), .outData_70(wire_con_in_stage1[70]), .outData_71(wire_con_in_stage1[71]), .outData_72(wire_con_in_stage1[72]), .outData_73(wire_con_in_stage1[73]), .outData_74(wire_con_in_stage1[74]), .outData_75(wire_con_in_stage1[75]), .outData_76(wire_con_in_stage1[76]), .outData_77(wire_con_in_stage1[77]), .outData_78(wire_con_in_stage1[78]), .outData_79(wire_con_in_stage1[79]), .outData_80(wire_con_in_stage1[80]), .outData_81(wire_con_in_stage1[81]), .outData_82(wire_con_in_stage1[82]), .outData_83(wire_con_in_stage1[83]), .outData_84(wire_con_in_stage1[84]), .outData_85(wire_con_in_stage1[85]), .outData_86(wire_con_in_stage1[86]), .outData_87(wire_con_in_stage1[87]), .outData_88(wire_con_in_stage1[88]), .outData_89(wire_con_in_stage1[89]), .outData_90(wire_con_in_stage1[90]), .outData_91(wire_con_in_stage1[91]), .outData_92(wire_con_in_stage1[92]), .outData_93(wire_con_in_stage1[93]), .outData_94(wire_con_in_stage1[94]), .outData_95(wire_con_in_stage1[95]), .outData_96(wire_con_in_stage1[96]), .outData_97(wire_con_in_stage1[97]), .outData_98(wire_con_in_stage1[98]), .outData_99(wire_con_in_stage1[99]), .outData_100(wire_con_in_stage1[100]), .outData_101(wire_con_in_stage1[101]), .outData_102(wire_con_in_stage1[102]), .outData_103(wire_con_in_stage1[103]), .outData_104(wire_con_in_stage1[104]), .outData_105(wire_con_in_stage1[105]), .outData_106(wire_con_in_stage1[106]), .outData_107(wire_con_in_stage1[107]), .outData_108(wire_con_in_stage1[108]), .outData_109(wire_con_in_stage1[109]), .outData_110(wire_con_in_stage1[110]), .outData_111(wire_con_in_stage1[111]), .outData_112(wire_con_in_stage1[112]), .outData_113(wire_con_in_stage1[113]), .outData_114(wire_con_in_stage1[114]), .outData_115(wire_con_in_stage1[115]), .outData_116(wire_con_in_stage1[116]), .outData_117(wire_con_in_stage1[117]), .outData_118(wire_con_in_stage1[118]), .outData_119(wire_con_in_stage1[119]), .outData_120(wire_con_in_stage1[120]), .outData_121(wire_con_in_stage1[121]), .outData_122(wire_con_in_stage1[122]), .outData_123(wire_con_in_stage1[123]), .outData_124(wire_con_in_stage1[124]), .outData_125(wire_con_in_stage1[125]), .outData_126(wire_con_in_stage1[126]), .outData_127(wire_con_in_stage1[127]), .outData_128(wire_con_in_stage1[128]), .outData_129(wire_con_in_stage1[129]), .outData_130(wire_con_in_stage1[130]), .outData_131(wire_con_in_stage1[131]), .outData_132(wire_con_in_stage1[132]), .outData_133(wire_con_in_stage1[133]), .outData_134(wire_con_in_stage1[134]), .outData_135(wire_con_in_stage1[135]), .outData_136(wire_con_in_stage1[136]), .outData_137(wire_con_in_stage1[137]), .outData_138(wire_con_in_stage1[138]), .outData_139(wire_con_in_stage1[139]), .outData_140(wire_con_in_stage1[140]), .outData_141(wire_con_in_stage1[141]), .outData_142(wire_con_in_stage1[142]), .outData_143(wire_con_in_stage1[143]), .outData_144(wire_con_in_stage1[144]), .outData_145(wire_con_in_stage1[145]), .outData_146(wire_con_in_stage1[146]), .outData_147(wire_con_in_stage1[147]), .outData_148(wire_con_in_stage1[148]), .outData_149(wire_con_in_stage1[149]), .outData_150(wire_con_in_stage1[150]), .outData_151(wire_con_in_stage1[151]), .outData_152(wire_con_in_stage1[152]), .outData_153(wire_con_in_stage1[153]), .outData_154(wire_con_in_stage1[154]), .outData_155(wire_con_in_stage1[155]), .outData_156(wire_con_in_stage1[156]), .outData_157(wire_con_in_stage1[157]), .outData_158(wire_con_in_stage1[158]), .outData_159(wire_con_in_stage1[159]), .outData_160(wire_con_in_stage1[160]), .outData_161(wire_con_in_stage1[161]), .outData_162(wire_con_in_stage1[162]), .outData_163(wire_con_in_stage1[163]), .outData_164(wire_con_in_stage1[164]), .outData_165(wire_con_in_stage1[165]), .outData_166(wire_con_in_stage1[166]), .outData_167(wire_con_in_stage1[167]), .outData_168(wire_con_in_stage1[168]), .outData_169(wire_con_in_stage1[169]), .outData_170(wire_con_in_stage1[170]), .outData_171(wire_con_in_stage1[171]), .outData_172(wire_con_in_stage1[172]), .outData_173(wire_con_in_stage1[173]), .outData_174(wire_con_in_stage1[174]), .outData_175(wire_con_in_stage1[175]), .outData_176(wire_con_in_stage1[176]), .outData_177(wire_con_in_stage1[177]), .outData_178(wire_con_in_stage1[178]), .outData_179(wire_con_in_stage1[179]), .outData_180(wire_con_in_stage1[180]), .outData_181(wire_con_in_stage1[181]), .outData_182(wire_con_in_stage1[182]), .outData_183(wire_con_in_stage1[183]), .outData_184(wire_con_in_stage1[184]), .outData_185(wire_con_in_stage1[185]), .outData_186(wire_con_in_stage1[186]), .outData_187(wire_con_in_stage1[187]), .outData_188(wire_con_in_stage1[188]), .outData_189(wire_con_in_stage1[189]), .outData_190(wire_con_in_stage1[190]), .outData_191(wire_con_in_stage1[191]), .outData_192(wire_con_in_stage1[192]), .outData_193(wire_con_in_stage1[193]), .outData_194(wire_con_in_stage1[194]), .outData_195(wire_con_in_stage1[195]), .outData_196(wire_con_in_stage1[196]), .outData_197(wire_con_in_stage1[197]), .outData_198(wire_con_in_stage1[198]), .outData_199(wire_con_in_stage1[199]), .outData_200(wire_con_in_stage1[200]), .outData_201(wire_con_in_stage1[201]), .outData_202(wire_con_in_stage1[202]), .outData_203(wire_con_in_stage1[203]), .outData_204(wire_con_in_stage1[204]), .outData_205(wire_con_in_stage1[205]), .outData_206(wire_con_in_stage1[206]), .outData_207(wire_con_in_stage1[207]), .outData_208(wire_con_in_stage1[208]), .outData_209(wire_con_in_stage1[209]), .outData_210(wire_con_in_stage1[210]), .outData_211(wire_con_in_stage1[211]), .outData_212(wire_con_in_stage1[212]), .outData_213(wire_con_in_stage1[213]), .outData_214(wire_con_in_stage1[214]), .outData_215(wire_con_in_stage1[215]), .outData_216(wire_con_in_stage1[216]), .outData_217(wire_con_in_stage1[217]), .outData_218(wire_con_in_stage1[218]), .outData_219(wire_con_in_stage1[219]), .outData_220(wire_con_in_stage1[220]), .outData_221(wire_con_in_stage1[221]), .outData_222(wire_con_in_stage1[222]), .outData_223(wire_con_in_stage1[223]), .outData_224(wire_con_in_stage1[224]), .outData_225(wire_con_in_stage1[225]), .outData_226(wire_con_in_stage1[226]), .outData_227(wire_con_in_stage1[227]), .outData_228(wire_con_in_stage1[228]), .outData_229(wire_con_in_stage1[229]), .outData_230(wire_con_in_stage1[230]), .outData_231(wire_con_in_stage1[231]), .outData_232(wire_con_in_stage1[232]), .outData_233(wire_con_in_stage1[233]), .outData_234(wire_con_in_stage1[234]), .outData_235(wire_con_in_stage1[235]), .outData_236(wire_con_in_stage1[236]), .outData_237(wire_con_in_stage1[237]), .outData_238(wire_con_in_stage1[238]), .outData_239(wire_con_in_stage1[239]), .outData_240(wire_con_in_stage1[240]), .outData_241(wire_con_in_stage1[241]), .outData_242(wire_con_in_stage1[242]), .outData_243(wire_con_in_stage1[243]), .outData_244(wire_con_in_stage1[244]), .outData_245(wire_con_in_stage1[245]), .outData_246(wire_con_in_stage1[246]), .outData_247(wire_con_in_stage1[247]), .outData_248(wire_con_in_stage1[248]), .outData_249(wire_con_in_stage1[249]), .outData_250(wire_con_in_stage1[250]), .outData_251(wire_con_in_stage1[251]), .outData_252(wire_con_in_stage1[252]), .outData_253(wire_con_in_stage1[253]), .outData_254(wire_con_in_stage1[254]), .outData_255(wire_con_in_stage1[255]), 
        .in_start(in_start_stage1), .out_start(con_in_start_stage1), .ctrl(wire_ctrl_stage1), .clk(clk), .rst(rst));
  
  wireCon_dp256_st1_L wire_stage_1(
        .inData_0(wire_con_in_stage1[0]), .inData_1(wire_con_in_stage1[1]), .inData_2(wire_con_in_stage1[2]), .inData_3(wire_con_in_stage1[3]), .inData_4(wire_con_in_stage1[4]), .inData_5(wire_con_in_stage1[5]), .inData_6(wire_con_in_stage1[6]), .inData_7(wire_con_in_stage1[7]), .inData_8(wire_con_in_stage1[8]), .inData_9(wire_con_in_stage1[9]), .inData_10(wire_con_in_stage1[10]), .inData_11(wire_con_in_stage1[11]), .inData_12(wire_con_in_stage1[12]), .inData_13(wire_con_in_stage1[13]), .inData_14(wire_con_in_stage1[14]), .inData_15(wire_con_in_stage1[15]), .inData_16(wire_con_in_stage1[16]), .inData_17(wire_con_in_stage1[17]), .inData_18(wire_con_in_stage1[18]), .inData_19(wire_con_in_stage1[19]), .inData_20(wire_con_in_stage1[20]), .inData_21(wire_con_in_stage1[21]), .inData_22(wire_con_in_stage1[22]), .inData_23(wire_con_in_stage1[23]), .inData_24(wire_con_in_stage1[24]), .inData_25(wire_con_in_stage1[25]), .inData_26(wire_con_in_stage1[26]), .inData_27(wire_con_in_stage1[27]), .inData_28(wire_con_in_stage1[28]), .inData_29(wire_con_in_stage1[29]), .inData_30(wire_con_in_stage1[30]), .inData_31(wire_con_in_stage1[31]), .inData_32(wire_con_in_stage1[32]), .inData_33(wire_con_in_stage1[33]), .inData_34(wire_con_in_stage1[34]), .inData_35(wire_con_in_stage1[35]), .inData_36(wire_con_in_stage1[36]), .inData_37(wire_con_in_stage1[37]), .inData_38(wire_con_in_stage1[38]), .inData_39(wire_con_in_stage1[39]), .inData_40(wire_con_in_stage1[40]), .inData_41(wire_con_in_stage1[41]), .inData_42(wire_con_in_stage1[42]), .inData_43(wire_con_in_stage1[43]), .inData_44(wire_con_in_stage1[44]), .inData_45(wire_con_in_stage1[45]), .inData_46(wire_con_in_stage1[46]), .inData_47(wire_con_in_stage1[47]), .inData_48(wire_con_in_stage1[48]), .inData_49(wire_con_in_stage1[49]), .inData_50(wire_con_in_stage1[50]), .inData_51(wire_con_in_stage1[51]), .inData_52(wire_con_in_stage1[52]), .inData_53(wire_con_in_stage1[53]), .inData_54(wire_con_in_stage1[54]), .inData_55(wire_con_in_stage1[55]), .inData_56(wire_con_in_stage1[56]), .inData_57(wire_con_in_stage1[57]), .inData_58(wire_con_in_stage1[58]), .inData_59(wire_con_in_stage1[59]), .inData_60(wire_con_in_stage1[60]), .inData_61(wire_con_in_stage1[61]), .inData_62(wire_con_in_stage1[62]), .inData_63(wire_con_in_stage1[63]), .inData_64(wire_con_in_stage1[64]), .inData_65(wire_con_in_stage1[65]), .inData_66(wire_con_in_stage1[66]), .inData_67(wire_con_in_stage1[67]), .inData_68(wire_con_in_stage1[68]), .inData_69(wire_con_in_stage1[69]), .inData_70(wire_con_in_stage1[70]), .inData_71(wire_con_in_stage1[71]), .inData_72(wire_con_in_stage1[72]), .inData_73(wire_con_in_stage1[73]), .inData_74(wire_con_in_stage1[74]), .inData_75(wire_con_in_stage1[75]), .inData_76(wire_con_in_stage1[76]), .inData_77(wire_con_in_stage1[77]), .inData_78(wire_con_in_stage1[78]), .inData_79(wire_con_in_stage1[79]), .inData_80(wire_con_in_stage1[80]), .inData_81(wire_con_in_stage1[81]), .inData_82(wire_con_in_stage1[82]), .inData_83(wire_con_in_stage1[83]), .inData_84(wire_con_in_stage1[84]), .inData_85(wire_con_in_stage1[85]), .inData_86(wire_con_in_stage1[86]), .inData_87(wire_con_in_stage1[87]), .inData_88(wire_con_in_stage1[88]), .inData_89(wire_con_in_stage1[89]), .inData_90(wire_con_in_stage1[90]), .inData_91(wire_con_in_stage1[91]), .inData_92(wire_con_in_stage1[92]), .inData_93(wire_con_in_stage1[93]), .inData_94(wire_con_in_stage1[94]), .inData_95(wire_con_in_stage1[95]), .inData_96(wire_con_in_stage1[96]), .inData_97(wire_con_in_stage1[97]), .inData_98(wire_con_in_stage1[98]), .inData_99(wire_con_in_stage1[99]), .inData_100(wire_con_in_stage1[100]), .inData_101(wire_con_in_stage1[101]), .inData_102(wire_con_in_stage1[102]), .inData_103(wire_con_in_stage1[103]), .inData_104(wire_con_in_stage1[104]), .inData_105(wire_con_in_stage1[105]), .inData_106(wire_con_in_stage1[106]), .inData_107(wire_con_in_stage1[107]), .inData_108(wire_con_in_stage1[108]), .inData_109(wire_con_in_stage1[109]), .inData_110(wire_con_in_stage1[110]), .inData_111(wire_con_in_stage1[111]), .inData_112(wire_con_in_stage1[112]), .inData_113(wire_con_in_stage1[113]), .inData_114(wire_con_in_stage1[114]), .inData_115(wire_con_in_stage1[115]), .inData_116(wire_con_in_stage1[116]), .inData_117(wire_con_in_stage1[117]), .inData_118(wire_con_in_stage1[118]), .inData_119(wire_con_in_stage1[119]), .inData_120(wire_con_in_stage1[120]), .inData_121(wire_con_in_stage1[121]), .inData_122(wire_con_in_stage1[122]), .inData_123(wire_con_in_stage1[123]), .inData_124(wire_con_in_stage1[124]), .inData_125(wire_con_in_stage1[125]), .inData_126(wire_con_in_stage1[126]), .inData_127(wire_con_in_stage1[127]), .inData_128(wire_con_in_stage1[128]), .inData_129(wire_con_in_stage1[129]), .inData_130(wire_con_in_stage1[130]), .inData_131(wire_con_in_stage1[131]), .inData_132(wire_con_in_stage1[132]), .inData_133(wire_con_in_stage1[133]), .inData_134(wire_con_in_stage1[134]), .inData_135(wire_con_in_stage1[135]), .inData_136(wire_con_in_stage1[136]), .inData_137(wire_con_in_stage1[137]), .inData_138(wire_con_in_stage1[138]), .inData_139(wire_con_in_stage1[139]), .inData_140(wire_con_in_stage1[140]), .inData_141(wire_con_in_stage1[141]), .inData_142(wire_con_in_stage1[142]), .inData_143(wire_con_in_stage1[143]), .inData_144(wire_con_in_stage1[144]), .inData_145(wire_con_in_stage1[145]), .inData_146(wire_con_in_stage1[146]), .inData_147(wire_con_in_stage1[147]), .inData_148(wire_con_in_stage1[148]), .inData_149(wire_con_in_stage1[149]), .inData_150(wire_con_in_stage1[150]), .inData_151(wire_con_in_stage1[151]), .inData_152(wire_con_in_stage1[152]), .inData_153(wire_con_in_stage1[153]), .inData_154(wire_con_in_stage1[154]), .inData_155(wire_con_in_stage1[155]), .inData_156(wire_con_in_stage1[156]), .inData_157(wire_con_in_stage1[157]), .inData_158(wire_con_in_stage1[158]), .inData_159(wire_con_in_stage1[159]), .inData_160(wire_con_in_stage1[160]), .inData_161(wire_con_in_stage1[161]), .inData_162(wire_con_in_stage1[162]), .inData_163(wire_con_in_stage1[163]), .inData_164(wire_con_in_stage1[164]), .inData_165(wire_con_in_stage1[165]), .inData_166(wire_con_in_stage1[166]), .inData_167(wire_con_in_stage1[167]), .inData_168(wire_con_in_stage1[168]), .inData_169(wire_con_in_stage1[169]), .inData_170(wire_con_in_stage1[170]), .inData_171(wire_con_in_stage1[171]), .inData_172(wire_con_in_stage1[172]), .inData_173(wire_con_in_stage1[173]), .inData_174(wire_con_in_stage1[174]), .inData_175(wire_con_in_stage1[175]), .inData_176(wire_con_in_stage1[176]), .inData_177(wire_con_in_stage1[177]), .inData_178(wire_con_in_stage1[178]), .inData_179(wire_con_in_stage1[179]), .inData_180(wire_con_in_stage1[180]), .inData_181(wire_con_in_stage1[181]), .inData_182(wire_con_in_stage1[182]), .inData_183(wire_con_in_stage1[183]), .inData_184(wire_con_in_stage1[184]), .inData_185(wire_con_in_stage1[185]), .inData_186(wire_con_in_stage1[186]), .inData_187(wire_con_in_stage1[187]), .inData_188(wire_con_in_stage1[188]), .inData_189(wire_con_in_stage1[189]), .inData_190(wire_con_in_stage1[190]), .inData_191(wire_con_in_stage1[191]), .inData_192(wire_con_in_stage1[192]), .inData_193(wire_con_in_stage1[193]), .inData_194(wire_con_in_stage1[194]), .inData_195(wire_con_in_stage1[195]), .inData_196(wire_con_in_stage1[196]), .inData_197(wire_con_in_stage1[197]), .inData_198(wire_con_in_stage1[198]), .inData_199(wire_con_in_stage1[199]), .inData_200(wire_con_in_stage1[200]), .inData_201(wire_con_in_stage1[201]), .inData_202(wire_con_in_stage1[202]), .inData_203(wire_con_in_stage1[203]), .inData_204(wire_con_in_stage1[204]), .inData_205(wire_con_in_stage1[205]), .inData_206(wire_con_in_stage1[206]), .inData_207(wire_con_in_stage1[207]), .inData_208(wire_con_in_stage1[208]), .inData_209(wire_con_in_stage1[209]), .inData_210(wire_con_in_stage1[210]), .inData_211(wire_con_in_stage1[211]), .inData_212(wire_con_in_stage1[212]), .inData_213(wire_con_in_stage1[213]), .inData_214(wire_con_in_stage1[214]), .inData_215(wire_con_in_stage1[215]), .inData_216(wire_con_in_stage1[216]), .inData_217(wire_con_in_stage1[217]), .inData_218(wire_con_in_stage1[218]), .inData_219(wire_con_in_stage1[219]), .inData_220(wire_con_in_stage1[220]), .inData_221(wire_con_in_stage1[221]), .inData_222(wire_con_in_stage1[222]), .inData_223(wire_con_in_stage1[223]), .inData_224(wire_con_in_stage1[224]), .inData_225(wire_con_in_stage1[225]), .inData_226(wire_con_in_stage1[226]), .inData_227(wire_con_in_stage1[227]), .inData_228(wire_con_in_stage1[228]), .inData_229(wire_con_in_stage1[229]), .inData_230(wire_con_in_stage1[230]), .inData_231(wire_con_in_stage1[231]), .inData_232(wire_con_in_stage1[232]), .inData_233(wire_con_in_stage1[233]), .inData_234(wire_con_in_stage1[234]), .inData_235(wire_con_in_stage1[235]), .inData_236(wire_con_in_stage1[236]), .inData_237(wire_con_in_stage1[237]), .inData_238(wire_con_in_stage1[238]), .inData_239(wire_con_in_stage1[239]), .inData_240(wire_con_in_stage1[240]), .inData_241(wire_con_in_stage1[241]), .inData_242(wire_con_in_stage1[242]), .inData_243(wire_con_in_stage1[243]), .inData_244(wire_con_in_stage1[244]), .inData_245(wire_con_in_stage1[245]), .inData_246(wire_con_in_stage1[246]), .inData_247(wire_con_in_stage1[247]), .inData_248(wire_con_in_stage1[248]), .inData_249(wire_con_in_stage1[249]), .inData_250(wire_con_in_stage1[250]), .inData_251(wire_con_in_stage1[251]), .inData_252(wire_con_in_stage1[252]), .inData_253(wire_con_in_stage1[253]), .inData_254(wire_con_in_stage1[254]), .inData_255(wire_con_in_stage1[255]), 
        .outData_0(wire_con_out_stage1[0]), .outData_1(wire_con_out_stage1[1]), .outData_2(wire_con_out_stage1[2]), .outData_3(wire_con_out_stage1[3]), .outData_4(wire_con_out_stage1[4]), .outData_5(wire_con_out_stage1[5]), .outData_6(wire_con_out_stage1[6]), .outData_7(wire_con_out_stage1[7]), .outData_8(wire_con_out_stage1[8]), .outData_9(wire_con_out_stage1[9]), .outData_10(wire_con_out_stage1[10]), .outData_11(wire_con_out_stage1[11]), .outData_12(wire_con_out_stage1[12]), .outData_13(wire_con_out_stage1[13]), .outData_14(wire_con_out_stage1[14]), .outData_15(wire_con_out_stage1[15]), .outData_16(wire_con_out_stage1[16]), .outData_17(wire_con_out_stage1[17]), .outData_18(wire_con_out_stage1[18]), .outData_19(wire_con_out_stage1[19]), .outData_20(wire_con_out_stage1[20]), .outData_21(wire_con_out_stage1[21]), .outData_22(wire_con_out_stage1[22]), .outData_23(wire_con_out_stage1[23]), .outData_24(wire_con_out_stage1[24]), .outData_25(wire_con_out_stage1[25]), .outData_26(wire_con_out_stage1[26]), .outData_27(wire_con_out_stage1[27]), .outData_28(wire_con_out_stage1[28]), .outData_29(wire_con_out_stage1[29]), .outData_30(wire_con_out_stage1[30]), .outData_31(wire_con_out_stage1[31]), .outData_32(wire_con_out_stage1[32]), .outData_33(wire_con_out_stage1[33]), .outData_34(wire_con_out_stage1[34]), .outData_35(wire_con_out_stage1[35]), .outData_36(wire_con_out_stage1[36]), .outData_37(wire_con_out_stage1[37]), .outData_38(wire_con_out_stage1[38]), .outData_39(wire_con_out_stage1[39]), .outData_40(wire_con_out_stage1[40]), .outData_41(wire_con_out_stage1[41]), .outData_42(wire_con_out_stage1[42]), .outData_43(wire_con_out_stage1[43]), .outData_44(wire_con_out_stage1[44]), .outData_45(wire_con_out_stage1[45]), .outData_46(wire_con_out_stage1[46]), .outData_47(wire_con_out_stage1[47]), .outData_48(wire_con_out_stage1[48]), .outData_49(wire_con_out_stage1[49]), .outData_50(wire_con_out_stage1[50]), .outData_51(wire_con_out_stage1[51]), .outData_52(wire_con_out_stage1[52]), .outData_53(wire_con_out_stage1[53]), .outData_54(wire_con_out_stage1[54]), .outData_55(wire_con_out_stage1[55]), .outData_56(wire_con_out_stage1[56]), .outData_57(wire_con_out_stage1[57]), .outData_58(wire_con_out_stage1[58]), .outData_59(wire_con_out_stage1[59]), .outData_60(wire_con_out_stage1[60]), .outData_61(wire_con_out_stage1[61]), .outData_62(wire_con_out_stage1[62]), .outData_63(wire_con_out_stage1[63]), .outData_64(wire_con_out_stage1[64]), .outData_65(wire_con_out_stage1[65]), .outData_66(wire_con_out_stage1[66]), .outData_67(wire_con_out_stage1[67]), .outData_68(wire_con_out_stage1[68]), .outData_69(wire_con_out_stage1[69]), .outData_70(wire_con_out_stage1[70]), .outData_71(wire_con_out_stage1[71]), .outData_72(wire_con_out_stage1[72]), .outData_73(wire_con_out_stage1[73]), .outData_74(wire_con_out_stage1[74]), .outData_75(wire_con_out_stage1[75]), .outData_76(wire_con_out_stage1[76]), .outData_77(wire_con_out_stage1[77]), .outData_78(wire_con_out_stage1[78]), .outData_79(wire_con_out_stage1[79]), .outData_80(wire_con_out_stage1[80]), .outData_81(wire_con_out_stage1[81]), .outData_82(wire_con_out_stage1[82]), .outData_83(wire_con_out_stage1[83]), .outData_84(wire_con_out_stage1[84]), .outData_85(wire_con_out_stage1[85]), .outData_86(wire_con_out_stage1[86]), .outData_87(wire_con_out_stage1[87]), .outData_88(wire_con_out_stage1[88]), .outData_89(wire_con_out_stage1[89]), .outData_90(wire_con_out_stage1[90]), .outData_91(wire_con_out_stage1[91]), .outData_92(wire_con_out_stage1[92]), .outData_93(wire_con_out_stage1[93]), .outData_94(wire_con_out_stage1[94]), .outData_95(wire_con_out_stage1[95]), .outData_96(wire_con_out_stage1[96]), .outData_97(wire_con_out_stage1[97]), .outData_98(wire_con_out_stage1[98]), .outData_99(wire_con_out_stage1[99]), .outData_100(wire_con_out_stage1[100]), .outData_101(wire_con_out_stage1[101]), .outData_102(wire_con_out_stage1[102]), .outData_103(wire_con_out_stage1[103]), .outData_104(wire_con_out_stage1[104]), .outData_105(wire_con_out_stage1[105]), .outData_106(wire_con_out_stage1[106]), .outData_107(wire_con_out_stage1[107]), .outData_108(wire_con_out_stage1[108]), .outData_109(wire_con_out_stage1[109]), .outData_110(wire_con_out_stage1[110]), .outData_111(wire_con_out_stage1[111]), .outData_112(wire_con_out_stage1[112]), .outData_113(wire_con_out_stage1[113]), .outData_114(wire_con_out_stage1[114]), .outData_115(wire_con_out_stage1[115]), .outData_116(wire_con_out_stage1[116]), .outData_117(wire_con_out_stage1[117]), .outData_118(wire_con_out_stage1[118]), .outData_119(wire_con_out_stage1[119]), .outData_120(wire_con_out_stage1[120]), .outData_121(wire_con_out_stage1[121]), .outData_122(wire_con_out_stage1[122]), .outData_123(wire_con_out_stage1[123]), .outData_124(wire_con_out_stage1[124]), .outData_125(wire_con_out_stage1[125]), .outData_126(wire_con_out_stage1[126]), .outData_127(wire_con_out_stage1[127]), .outData_128(wire_con_out_stage1[128]), .outData_129(wire_con_out_stage1[129]), .outData_130(wire_con_out_stage1[130]), .outData_131(wire_con_out_stage1[131]), .outData_132(wire_con_out_stage1[132]), .outData_133(wire_con_out_stage1[133]), .outData_134(wire_con_out_stage1[134]), .outData_135(wire_con_out_stage1[135]), .outData_136(wire_con_out_stage1[136]), .outData_137(wire_con_out_stage1[137]), .outData_138(wire_con_out_stage1[138]), .outData_139(wire_con_out_stage1[139]), .outData_140(wire_con_out_stage1[140]), .outData_141(wire_con_out_stage1[141]), .outData_142(wire_con_out_stage1[142]), .outData_143(wire_con_out_stage1[143]), .outData_144(wire_con_out_stage1[144]), .outData_145(wire_con_out_stage1[145]), .outData_146(wire_con_out_stage1[146]), .outData_147(wire_con_out_stage1[147]), .outData_148(wire_con_out_stage1[148]), .outData_149(wire_con_out_stage1[149]), .outData_150(wire_con_out_stage1[150]), .outData_151(wire_con_out_stage1[151]), .outData_152(wire_con_out_stage1[152]), .outData_153(wire_con_out_stage1[153]), .outData_154(wire_con_out_stage1[154]), .outData_155(wire_con_out_stage1[155]), .outData_156(wire_con_out_stage1[156]), .outData_157(wire_con_out_stage1[157]), .outData_158(wire_con_out_stage1[158]), .outData_159(wire_con_out_stage1[159]), .outData_160(wire_con_out_stage1[160]), .outData_161(wire_con_out_stage1[161]), .outData_162(wire_con_out_stage1[162]), .outData_163(wire_con_out_stage1[163]), .outData_164(wire_con_out_stage1[164]), .outData_165(wire_con_out_stage1[165]), .outData_166(wire_con_out_stage1[166]), .outData_167(wire_con_out_stage1[167]), .outData_168(wire_con_out_stage1[168]), .outData_169(wire_con_out_stage1[169]), .outData_170(wire_con_out_stage1[170]), .outData_171(wire_con_out_stage1[171]), .outData_172(wire_con_out_stage1[172]), .outData_173(wire_con_out_stage1[173]), .outData_174(wire_con_out_stage1[174]), .outData_175(wire_con_out_stage1[175]), .outData_176(wire_con_out_stage1[176]), .outData_177(wire_con_out_stage1[177]), .outData_178(wire_con_out_stage1[178]), .outData_179(wire_con_out_stage1[179]), .outData_180(wire_con_out_stage1[180]), .outData_181(wire_con_out_stage1[181]), .outData_182(wire_con_out_stage1[182]), .outData_183(wire_con_out_stage1[183]), .outData_184(wire_con_out_stage1[184]), .outData_185(wire_con_out_stage1[185]), .outData_186(wire_con_out_stage1[186]), .outData_187(wire_con_out_stage1[187]), .outData_188(wire_con_out_stage1[188]), .outData_189(wire_con_out_stage1[189]), .outData_190(wire_con_out_stage1[190]), .outData_191(wire_con_out_stage1[191]), .outData_192(wire_con_out_stage1[192]), .outData_193(wire_con_out_stage1[193]), .outData_194(wire_con_out_stage1[194]), .outData_195(wire_con_out_stage1[195]), .outData_196(wire_con_out_stage1[196]), .outData_197(wire_con_out_stage1[197]), .outData_198(wire_con_out_stage1[198]), .outData_199(wire_con_out_stage1[199]), .outData_200(wire_con_out_stage1[200]), .outData_201(wire_con_out_stage1[201]), .outData_202(wire_con_out_stage1[202]), .outData_203(wire_con_out_stage1[203]), .outData_204(wire_con_out_stage1[204]), .outData_205(wire_con_out_stage1[205]), .outData_206(wire_con_out_stage1[206]), .outData_207(wire_con_out_stage1[207]), .outData_208(wire_con_out_stage1[208]), .outData_209(wire_con_out_stage1[209]), .outData_210(wire_con_out_stage1[210]), .outData_211(wire_con_out_stage1[211]), .outData_212(wire_con_out_stage1[212]), .outData_213(wire_con_out_stage1[213]), .outData_214(wire_con_out_stage1[214]), .outData_215(wire_con_out_stage1[215]), .outData_216(wire_con_out_stage1[216]), .outData_217(wire_con_out_stage1[217]), .outData_218(wire_con_out_stage1[218]), .outData_219(wire_con_out_stage1[219]), .outData_220(wire_con_out_stage1[220]), .outData_221(wire_con_out_stage1[221]), .outData_222(wire_con_out_stage1[222]), .outData_223(wire_con_out_stage1[223]), .outData_224(wire_con_out_stage1[224]), .outData_225(wire_con_out_stage1[225]), .outData_226(wire_con_out_stage1[226]), .outData_227(wire_con_out_stage1[227]), .outData_228(wire_con_out_stage1[228]), .outData_229(wire_con_out_stage1[229]), .outData_230(wire_con_out_stage1[230]), .outData_231(wire_con_out_stage1[231]), .outData_232(wire_con_out_stage1[232]), .outData_233(wire_con_out_stage1[233]), .outData_234(wire_con_out_stage1[234]), .outData_235(wire_con_out_stage1[235]), .outData_236(wire_con_out_stage1[236]), .outData_237(wire_con_out_stage1[237]), .outData_238(wire_con_out_stage1[238]), .outData_239(wire_con_out_stage1[239]), .outData_240(wire_con_out_stage1[240]), .outData_241(wire_con_out_stage1[241]), .outData_242(wire_con_out_stage1[242]), .outData_243(wire_con_out_stage1[243]), .outData_244(wire_con_out_stage1[244]), .outData_245(wire_con_out_stage1[245]), .outData_246(wire_con_out_stage1[246]), .outData_247(wire_con_out_stage1[247]), .outData_248(wire_con_out_stage1[248]), .outData_249(wire_con_out_stage1[249]), .outData_250(wire_con_out_stage1[250]), .outData_251(wire_con_out_stage1[251]), .outData_252(wire_con_out_stage1[252]), .outData_253(wire_con_out_stage1[253]), .outData_254(wire_con_out_stage1[254]), .outData_255(wire_con_out_stage1[255]), 
        .in_start(con_in_start_stage1), .out_start(in_start_stage2), .clk(clk), .rst(rst)); 

  
  assign wire_ctrl_stage1[0] = counter_w[6]; 
  assign wire_ctrl_stage1[1] = counter_w[6]; 
  assign wire_ctrl_stage1[2] = counter_w[6]; 
  assign wire_ctrl_stage1[3] = counter_w[6]; 
  assign wire_ctrl_stage1[4] = counter_w[6]; 
  assign wire_ctrl_stage1[5] = counter_w[6]; 
  assign wire_ctrl_stage1[6] = counter_w[6]; 
  assign wire_ctrl_stage1[7] = counter_w[6]; 
  assign wire_ctrl_stage1[8] = counter_w[6]; 
  assign wire_ctrl_stage1[9] = counter_w[6]; 
  assign wire_ctrl_stage1[10] = counter_w[6]; 
  assign wire_ctrl_stage1[11] = counter_w[6]; 
  assign wire_ctrl_stage1[12] = counter_w[6]; 
  assign wire_ctrl_stage1[13] = counter_w[6]; 
  assign wire_ctrl_stage1[14] = counter_w[6]; 
  assign wire_ctrl_stage1[15] = counter_w[6]; 
  assign wire_ctrl_stage1[16] = counter_w[6]; 
  assign wire_ctrl_stage1[17] = counter_w[6]; 
  assign wire_ctrl_stage1[18] = counter_w[6]; 
  assign wire_ctrl_stage1[19] = counter_w[6]; 
  assign wire_ctrl_stage1[20] = counter_w[6]; 
  assign wire_ctrl_stage1[21] = counter_w[6]; 
  assign wire_ctrl_stage1[22] = counter_w[6]; 
  assign wire_ctrl_stage1[23] = counter_w[6]; 
  assign wire_ctrl_stage1[24] = counter_w[6]; 
  assign wire_ctrl_stage1[25] = counter_w[6]; 
  assign wire_ctrl_stage1[26] = counter_w[6]; 
  assign wire_ctrl_stage1[27] = counter_w[6]; 
  assign wire_ctrl_stage1[28] = counter_w[6]; 
  assign wire_ctrl_stage1[29] = counter_w[6]; 
  assign wire_ctrl_stage1[30] = counter_w[6]; 
  assign wire_ctrl_stage1[31] = counter_w[6]; 
  assign wire_ctrl_stage1[32] = counter_w[6]; 
  assign wire_ctrl_stage1[33] = counter_w[6]; 
  assign wire_ctrl_stage1[34] = counter_w[6]; 
  assign wire_ctrl_stage1[35] = counter_w[6]; 
  assign wire_ctrl_stage1[36] = counter_w[6]; 
  assign wire_ctrl_stage1[37] = counter_w[6]; 
  assign wire_ctrl_stage1[38] = counter_w[6]; 
  assign wire_ctrl_stage1[39] = counter_w[6]; 
  assign wire_ctrl_stage1[40] = counter_w[6]; 
  assign wire_ctrl_stage1[41] = counter_w[6]; 
  assign wire_ctrl_stage1[42] = counter_w[6]; 
  assign wire_ctrl_stage1[43] = counter_w[6]; 
  assign wire_ctrl_stage1[44] = counter_w[6]; 
  assign wire_ctrl_stage1[45] = counter_w[6]; 
  assign wire_ctrl_stage1[46] = counter_w[6]; 
  assign wire_ctrl_stage1[47] = counter_w[6]; 
  assign wire_ctrl_stage1[48] = counter_w[6]; 
  assign wire_ctrl_stage1[49] = counter_w[6]; 
  assign wire_ctrl_stage1[50] = counter_w[6]; 
  assign wire_ctrl_stage1[51] = counter_w[6]; 
  assign wire_ctrl_stage1[52] = counter_w[6]; 
  assign wire_ctrl_stage1[53] = counter_w[6]; 
  assign wire_ctrl_stage1[54] = counter_w[6]; 
  assign wire_ctrl_stage1[55] = counter_w[6]; 
  assign wire_ctrl_stage1[56] = counter_w[6]; 
  assign wire_ctrl_stage1[57] = counter_w[6]; 
  assign wire_ctrl_stage1[58] = counter_w[6]; 
  assign wire_ctrl_stage1[59] = counter_w[6]; 
  assign wire_ctrl_stage1[60] = counter_w[6]; 
  assign wire_ctrl_stage1[61] = counter_w[6]; 
  assign wire_ctrl_stage1[62] = counter_w[6]; 
  assign wire_ctrl_stage1[63] = counter_w[6]; 
  assign wire_ctrl_stage1[64] = counter_w[6]; 
  assign wire_ctrl_stage1[65] = counter_w[6]; 
  assign wire_ctrl_stage1[66] = counter_w[6]; 
  assign wire_ctrl_stage1[67] = counter_w[6]; 
  assign wire_ctrl_stage1[68] = counter_w[6]; 
  assign wire_ctrl_stage1[69] = counter_w[6]; 
  assign wire_ctrl_stage1[70] = counter_w[6]; 
  assign wire_ctrl_stage1[71] = counter_w[6]; 
  assign wire_ctrl_stage1[72] = counter_w[6]; 
  assign wire_ctrl_stage1[73] = counter_w[6]; 
  assign wire_ctrl_stage1[74] = counter_w[6]; 
  assign wire_ctrl_stage1[75] = counter_w[6]; 
  assign wire_ctrl_stage1[76] = counter_w[6]; 
  assign wire_ctrl_stage1[77] = counter_w[6]; 
  assign wire_ctrl_stage1[78] = counter_w[6]; 
  assign wire_ctrl_stage1[79] = counter_w[6]; 
  assign wire_ctrl_stage1[80] = counter_w[6]; 
  assign wire_ctrl_stage1[81] = counter_w[6]; 
  assign wire_ctrl_stage1[82] = counter_w[6]; 
  assign wire_ctrl_stage1[83] = counter_w[6]; 
  assign wire_ctrl_stage1[84] = counter_w[6]; 
  assign wire_ctrl_stage1[85] = counter_w[6]; 
  assign wire_ctrl_stage1[86] = counter_w[6]; 
  assign wire_ctrl_stage1[87] = counter_w[6]; 
  assign wire_ctrl_stage1[88] = counter_w[6]; 
  assign wire_ctrl_stage1[89] = counter_w[6]; 
  assign wire_ctrl_stage1[90] = counter_w[6]; 
  assign wire_ctrl_stage1[91] = counter_w[6]; 
  assign wire_ctrl_stage1[92] = counter_w[6]; 
  assign wire_ctrl_stage1[93] = counter_w[6]; 
  assign wire_ctrl_stage1[94] = counter_w[6]; 
  assign wire_ctrl_stage1[95] = counter_w[6]; 
  assign wire_ctrl_stage1[96] = counter_w[6]; 
  assign wire_ctrl_stage1[97] = counter_w[6]; 
  assign wire_ctrl_stage1[98] = counter_w[6]; 
  assign wire_ctrl_stage1[99] = counter_w[6]; 
  assign wire_ctrl_stage1[100] = counter_w[6]; 
  assign wire_ctrl_stage1[101] = counter_w[6]; 
  assign wire_ctrl_stage1[102] = counter_w[6]; 
  assign wire_ctrl_stage1[103] = counter_w[6]; 
  assign wire_ctrl_stage1[104] = counter_w[6]; 
  assign wire_ctrl_stage1[105] = counter_w[6]; 
  assign wire_ctrl_stage1[106] = counter_w[6]; 
  assign wire_ctrl_stage1[107] = counter_w[6]; 
  assign wire_ctrl_stage1[108] = counter_w[6]; 
  assign wire_ctrl_stage1[109] = counter_w[6]; 
  assign wire_ctrl_stage1[110] = counter_w[6]; 
  assign wire_ctrl_stage1[111] = counter_w[6]; 
  assign wire_ctrl_stage1[112] = counter_w[6]; 
  assign wire_ctrl_stage1[113] = counter_w[6]; 
  assign wire_ctrl_stage1[114] = counter_w[6]; 
  assign wire_ctrl_stage1[115] = counter_w[6]; 
  assign wire_ctrl_stage1[116] = counter_w[6]; 
  assign wire_ctrl_stage1[117] = counter_w[6]; 
  assign wire_ctrl_stage1[118] = counter_w[6]; 
  assign wire_ctrl_stage1[119] = counter_w[6]; 
  assign wire_ctrl_stage1[120] = counter_w[6]; 
  assign wire_ctrl_stage1[121] = counter_w[6]; 
  assign wire_ctrl_stage1[122] = counter_w[6]; 
  assign wire_ctrl_stage1[123] = counter_w[6]; 
  assign wire_ctrl_stage1[124] = counter_w[6]; 
  assign wire_ctrl_stage1[125] = counter_w[6]; 
  assign wire_ctrl_stage1[126] = counter_w[6]; 
  assign wire_ctrl_stage1[127] = counter_w[6]; 
  wire [DATA_WIDTH-1:0] wire_con_in_stage2[255:0];
  wire [DATA_WIDTH-1:0] wire_con_out_stage2[255:0];
  wire [127:0] wire_ctrl_stage2;

  switches_stage_st2_0_L switch_stage_2(
        .inData_0(wire_con_out_stage1[0]), .inData_1(wire_con_out_stage1[1]), .inData_2(wire_con_out_stage1[2]), .inData_3(wire_con_out_stage1[3]), .inData_4(wire_con_out_stage1[4]), .inData_5(wire_con_out_stage1[5]), .inData_6(wire_con_out_stage1[6]), .inData_7(wire_con_out_stage1[7]), .inData_8(wire_con_out_stage1[8]), .inData_9(wire_con_out_stage1[9]), .inData_10(wire_con_out_stage1[10]), .inData_11(wire_con_out_stage1[11]), .inData_12(wire_con_out_stage1[12]), .inData_13(wire_con_out_stage1[13]), .inData_14(wire_con_out_stage1[14]), .inData_15(wire_con_out_stage1[15]), .inData_16(wire_con_out_stage1[16]), .inData_17(wire_con_out_stage1[17]), .inData_18(wire_con_out_stage1[18]), .inData_19(wire_con_out_stage1[19]), .inData_20(wire_con_out_stage1[20]), .inData_21(wire_con_out_stage1[21]), .inData_22(wire_con_out_stage1[22]), .inData_23(wire_con_out_stage1[23]), .inData_24(wire_con_out_stage1[24]), .inData_25(wire_con_out_stage1[25]), .inData_26(wire_con_out_stage1[26]), .inData_27(wire_con_out_stage1[27]), .inData_28(wire_con_out_stage1[28]), .inData_29(wire_con_out_stage1[29]), .inData_30(wire_con_out_stage1[30]), .inData_31(wire_con_out_stage1[31]), .inData_32(wire_con_out_stage1[32]), .inData_33(wire_con_out_stage1[33]), .inData_34(wire_con_out_stage1[34]), .inData_35(wire_con_out_stage1[35]), .inData_36(wire_con_out_stage1[36]), .inData_37(wire_con_out_stage1[37]), .inData_38(wire_con_out_stage1[38]), .inData_39(wire_con_out_stage1[39]), .inData_40(wire_con_out_stage1[40]), .inData_41(wire_con_out_stage1[41]), .inData_42(wire_con_out_stage1[42]), .inData_43(wire_con_out_stage1[43]), .inData_44(wire_con_out_stage1[44]), .inData_45(wire_con_out_stage1[45]), .inData_46(wire_con_out_stage1[46]), .inData_47(wire_con_out_stage1[47]), .inData_48(wire_con_out_stage1[48]), .inData_49(wire_con_out_stage1[49]), .inData_50(wire_con_out_stage1[50]), .inData_51(wire_con_out_stage1[51]), .inData_52(wire_con_out_stage1[52]), .inData_53(wire_con_out_stage1[53]), .inData_54(wire_con_out_stage1[54]), .inData_55(wire_con_out_stage1[55]), .inData_56(wire_con_out_stage1[56]), .inData_57(wire_con_out_stage1[57]), .inData_58(wire_con_out_stage1[58]), .inData_59(wire_con_out_stage1[59]), .inData_60(wire_con_out_stage1[60]), .inData_61(wire_con_out_stage1[61]), .inData_62(wire_con_out_stage1[62]), .inData_63(wire_con_out_stage1[63]), .inData_64(wire_con_out_stage1[64]), .inData_65(wire_con_out_stage1[65]), .inData_66(wire_con_out_stage1[66]), .inData_67(wire_con_out_stage1[67]), .inData_68(wire_con_out_stage1[68]), .inData_69(wire_con_out_stage1[69]), .inData_70(wire_con_out_stage1[70]), .inData_71(wire_con_out_stage1[71]), .inData_72(wire_con_out_stage1[72]), .inData_73(wire_con_out_stage1[73]), .inData_74(wire_con_out_stage1[74]), .inData_75(wire_con_out_stage1[75]), .inData_76(wire_con_out_stage1[76]), .inData_77(wire_con_out_stage1[77]), .inData_78(wire_con_out_stage1[78]), .inData_79(wire_con_out_stage1[79]), .inData_80(wire_con_out_stage1[80]), .inData_81(wire_con_out_stage1[81]), .inData_82(wire_con_out_stage1[82]), .inData_83(wire_con_out_stage1[83]), .inData_84(wire_con_out_stage1[84]), .inData_85(wire_con_out_stage1[85]), .inData_86(wire_con_out_stage1[86]), .inData_87(wire_con_out_stage1[87]), .inData_88(wire_con_out_stage1[88]), .inData_89(wire_con_out_stage1[89]), .inData_90(wire_con_out_stage1[90]), .inData_91(wire_con_out_stage1[91]), .inData_92(wire_con_out_stage1[92]), .inData_93(wire_con_out_stage1[93]), .inData_94(wire_con_out_stage1[94]), .inData_95(wire_con_out_stage1[95]), .inData_96(wire_con_out_stage1[96]), .inData_97(wire_con_out_stage1[97]), .inData_98(wire_con_out_stage1[98]), .inData_99(wire_con_out_stage1[99]), .inData_100(wire_con_out_stage1[100]), .inData_101(wire_con_out_stage1[101]), .inData_102(wire_con_out_stage1[102]), .inData_103(wire_con_out_stage1[103]), .inData_104(wire_con_out_stage1[104]), .inData_105(wire_con_out_stage1[105]), .inData_106(wire_con_out_stage1[106]), .inData_107(wire_con_out_stage1[107]), .inData_108(wire_con_out_stage1[108]), .inData_109(wire_con_out_stage1[109]), .inData_110(wire_con_out_stage1[110]), .inData_111(wire_con_out_stage1[111]), .inData_112(wire_con_out_stage1[112]), .inData_113(wire_con_out_stage1[113]), .inData_114(wire_con_out_stage1[114]), .inData_115(wire_con_out_stage1[115]), .inData_116(wire_con_out_stage1[116]), .inData_117(wire_con_out_stage1[117]), .inData_118(wire_con_out_stage1[118]), .inData_119(wire_con_out_stage1[119]), .inData_120(wire_con_out_stage1[120]), .inData_121(wire_con_out_stage1[121]), .inData_122(wire_con_out_stage1[122]), .inData_123(wire_con_out_stage1[123]), .inData_124(wire_con_out_stage1[124]), .inData_125(wire_con_out_stage1[125]), .inData_126(wire_con_out_stage1[126]), .inData_127(wire_con_out_stage1[127]), .inData_128(wire_con_out_stage1[128]), .inData_129(wire_con_out_stage1[129]), .inData_130(wire_con_out_stage1[130]), .inData_131(wire_con_out_stage1[131]), .inData_132(wire_con_out_stage1[132]), .inData_133(wire_con_out_stage1[133]), .inData_134(wire_con_out_stage1[134]), .inData_135(wire_con_out_stage1[135]), .inData_136(wire_con_out_stage1[136]), .inData_137(wire_con_out_stage1[137]), .inData_138(wire_con_out_stage1[138]), .inData_139(wire_con_out_stage1[139]), .inData_140(wire_con_out_stage1[140]), .inData_141(wire_con_out_stage1[141]), .inData_142(wire_con_out_stage1[142]), .inData_143(wire_con_out_stage1[143]), .inData_144(wire_con_out_stage1[144]), .inData_145(wire_con_out_stage1[145]), .inData_146(wire_con_out_stage1[146]), .inData_147(wire_con_out_stage1[147]), .inData_148(wire_con_out_stage1[148]), .inData_149(wire_con_out_stage1[149]), .inData_150(wire_con_out_stage1[150]), .inData_151(wire_con_out_stage1[151]), .inData_152(wire_con_out_stage1[152]), .inData_153(wire_con_out_stage1[153]), .inData_154(wire_con_out_stage1[154]), .inData_155(wire_con_out_stage1[155]), .inData_156(wire_con_out_stage1[156]), .inData_157(wire_con_out_stage1[157]), .inData_158(wire_con_out_stage1[158]), .inData_159(wire_con_out_stage1[159]), .inData_160(wire_con_out_stage1[160]), .inData_161(wire_con_out_stage1[161]), .inData_162(wire_con_out_stage1[162]), .inData_163(wire_con_out_stage1[163]), .inData_164(wire_con_out_stage1[164]), .inData_165(wire_con_out_stage1[165]), .inData_166(wire_con_out_stage1[166]), .inData_167(wire_con_out_stage1[167]), .inData_168(wire_con_out_stage1[168]), .inData_169(wire_con_out_stage1[169]), .inData_170(wire_con_out_stage1[170]), .inData_171(wire_con_out_stage1[171]), .inData_172(wire_con_out_stage1[172]), .inData_173(wire_con_out_stage1[173]), .inData_174(wire_con_out_stage1[174]), .inData_175(wire_con_out_stage1[175]), .inData_176(wire_con_out_stage1[176]), .inData_177(wire_con_out_stage1[177]), .inData_178(wire_con_out_stage1[178]), .inData_179(wire_con_out_stage1[179]), .inData_180(wire_con_out_stage1[180]), .inData_181(wire_con_out_stage1[181]), .inData_182(wire_con_out_stage1[182]), .inData_183(wire_con_out_stage1[183]), .inData_184(wire_con_out_stage1[184]), .inData_185(wire_con_out_stage1[185]), .inData_186(wire_con_out_stage1[186]), .inData_187(wire_con_out_stage1[187]), .inData_188(wire_con_out_stage1[188]), .inData_189(wire_con_out_stage1[189]), .inData_190(wire_con_out_stage1[190]), .inData_191(wire_con_out_stage1[191]), .inData_192(wire_con_out_stage1[192]), .inData_193(wire_con_out_stage1[193]), .inData_194(wire_con_out_stage1[194]), .inData_195(wire_con_out_stage1[195]), .inData_196(wire_con_out_stage1[196]), .inData_197(wire_con_out_stage1[197]), .inData_198(wire_con_out_stage1[198]), .inData_199(wire_con_out_stage1[199]), .inData_200(wire_con_out_stage1[200]), .inData_201(wire_con_out_stage1[201]), .inData_202(wire_con_out_stage1[202]), .inData_203(wire_con_out_stage1[203]), .inData_204(wire_con_out_stage1[204]), .inData_205(wire_con_out_stage1[205]), .inData_206(wire_con_out_stage1[206]), .inData_207(wire_con_out_stage1[207]), .inData_208(wire_con_out_stage1[208]), .inData_209(wire_con_out_stage1[209]), .inData_210(wire_con_out_stage1[210]), .inData_211(wire_con_out_stage1[211]), .inData_212(wire_con_out_stage1[212]), .inData_213(wire_con_out_stage1[213]), .inData_214(wire_con_out_stage1[214]), .inData_215(wire_con_out_stage1[215]), .inData_216(wire_con_out_stage1[216]), .inData_217(wire_con_out_stage1[217]), .inData_218(wire_con_out_stage1[218]), .inData_219(wire_con_out_stage1[219]), .inData_220(wire_con_out_stage1[220]), .inData_221(wire_con_out_stage1[221]), .inData_222(wire_con_out_stage1[222]), .inData_223(wire_con_out_stage1[223]), .inData_224(wire_con_out_stage1[224]), .inData_225(wire_con_out_stage1[225]), .inData_226(wire_con_out_stage1[226]), .inData_227(wire_con_out_stage1[227]), .inData_228(wire_con_out_stage1[228]), .inData_229(wire_con_out_stage1[229]), .inData_230(wire_con_out_stage1[230]), .inData_231(wire_con_out_stage1[231]), .inData_232(wire_con_out_stage1[232]), .inData_233(wire_con_out_stage1[233]), .inData_234(wire_con_out_stage1[234]), .inData_235(wire_con_out_stage1[235]), .inData_236(wire_con_out_stage1[236]), .inData_237(wire_con_out_stage1[237]), .inData_238(wire_con_out_stage1[238]), .inData_239(wire_con_out_stage1[239]), .inData_240(wire_con_out_stage1[240]), .inData_241(wire_con_out_stage1[241]), .inData_242(wire_con_out_stage1[242]), .inData_243(wire_con_out_stage1[243]), .inData_244(wire_con_out_stage1[244]), .inData_245(wire_con_out_stage1[245]), .inData_246(wire_con_out_stage1[246]), .inData_247(wire_con_out_stage1[247]), .inData_248(wire_con_out_stage1[248]), .inData_249(wire_con_out_stage1[249]), .inData_250(wire_con_out_stage1[250]), .inData_251(wire_con_out_stage1[251]), .inData_252(wire_con_out_stage1[252]), .inData_253(wire_con_out_stage1[253]), .inData_254(wire_con_out_stage1[254]), .inData_255(wire_con_out_stage1[255]), 
        .outData_0(wire_con_in_stage2[0]), .outData_1(wire_con_in_stage2[1]), .outData_2(wire_con_in_stage2[2]), .outData_3(wire_con_in_stage2[3]), .outData_4(wire_con_in_stage2[4]), .outData_5(wire_con_in_stage2[5]), .outData_6(wire_con_in_stage2[6]), .outData_7(wire_con_in_stage2[7]), .outData_8(wire_con_in_stage2[8]), .outData_9(wire_con_in_stage2[9]), .outData_10(wire_con_in_stage2[10]), .outData_11(wire_con_in_stage2[11]), .outData_12(wire_con_in_stage2[12]), .outData_13(wire_con_in_stage2[13]), .outData_14(wire_con_in_stage2[14]), .outData_15(wire_con_in_stage2[15]), .outData_16(wire_con_in_stage2[16]), .outData_17(wire_con_in_stage2[17]), .outData_18(wire_con_in_stage2[18]), .outData_19(wire_con_in_stage2[19]), .outData_20(wire_con_in_stage2[20]), .outData_21(wire_con_in_stage2[21]), .outData_22(wire_con_in_stage2[22]), .outData_23(wire_con_in_stage2[23]), .outData_24(wire_con_in_stage2[24]), .outData_25(wire_con_in_stage2[25]), .outData_26(wire_con_in_stage2[26]), .outData_27(wire_con_in_stage2[27]), .outData_28(wire_con_in_stage2[28]), .outData_29(wire_con_in_stage2[29]), .outData_30(wire_con_in_stage2[30]), .outData_31(wire_con_in_stage2[31]), .outData_32(wire_con_in_stage2[32]), .outData_33(wire_con_in_stage2[33]), .outData_34(wire_con_in_stage2[34]), .outData_35(wire_con_in_stage2[35]), .outData_36(wire_con_in_stage2[36]), .outData_37(wire_con_in_stage2[37]), .outData_38(wire_con_in_stage2[38]), .outData_39(wire_con_in_stage2[39]), .outData_40(wire_con_in_stage2[40]), .outData_41(wire_con_in_stage2[41]), .outData_42(wire_con_in_stage2[42]), .outData_43(wire_con_in_stage2[43]), .outData_44(wire_con_in_stage2[44]), .outData_45(wire_con_in_stage2[45]), .outData_46(wire_con_in_stage2[46]), .outData_47(wire_con_in_stage2[47]), .outData_48(wire_con_in_stage2[48]), .outData_49(wire_con_in_stage2[49]), .outData_50(wire_con_in_stage2[50]), .outData_51(wire_con_in_stage2[51]), .outData_52(wire_con_in_stage2[52]), .outData_53(wire_con_in_stage2[53]), .outData_54(wire_con_in_stage2[54]), .outData_55(wire_con_in_stage2[55]), .outData_56(wire_con_in_stage2[56]), .outData_57(wire_con_in_stage2[57]), .outData_58(wire_con_in_stage2[58]), .outData_59(wire_con_in_stage2[59]), .outData_60(wire_con_in_stage2[60]), .outData_61(wire_con_in_stage2[61]), .outData_62(wire_con_in_stage2[62]), .outData_63(wire_con_in_stage2[63]), .outData_64(wire_con_in_stage2[64]), .outData_65(wire_con_in_stage2[65]), .outData_66(wire_con_in_stage2[66]), .outData_67(wire_con_in_stage2[67]), .outData_68(wire_con_in_stage2[68]), .outData_69(wire_con_in_stage2[69]), .outData_70(wire_con_in_stage2[70]), .outData_71(wire_con_in_stage2[71]), .outData_72(wire_con_in_stage2[72]), .outData_73(wire_con_in_stage2[73]), .outData_74(wire_con_in_stage2[74]), .outData_75(wire_con_in_stage2[75]), .outData_76(wire_con_in_stage2[76]), .outData_77(wire_con_in_stage2[77]), .outData_78(wire_con_in_stage2[78]), .outData_79(wire_con_in_stage2[79]), .outData_80(wire_con_in_stage2[80]), .outData_81(wire_con_in_stage2[81]), .outData_82(wire_con_in_stage2[82]), .outData_83(wire_con_in_stage2[83]), .outData_84(wire_con_in_stage2[84]), .outData_85(wire_con_in_stage2[85]), .outData_86(wire_con_in_stage2[86]), .outData_87(wire_con_in_stage2[87]), .outData_88(wire_con_in_stage2[88]), .outData_89(wire_con_in_stage2[89]), .outData_90(wire_con_in_stage2[90]), .outData_91(wire_con_in_stage2[91]), .outData_92(wire_con_in_stage2[92]), .outData_93(wire_con_in_stage2[93]), .outData_94(wire_con_in_stage2[94]), .outData_95(wire_con_in_stage2[95]), .outData_96(wire_con_in_stage2[96]), .outData_97(wire_con_in_stage2[97]), .outData_98(wire_con_in_stage2[98]), .outData_99(wire_con_in_stage2[99]), .outData_100(wire_con_in_stage2[100]), .outData_101(wire_con_in_stage2[101]), .outData_102(wire_con_in_stage2[102]), .outData_103(wire_con_in_stage2[103]), .outData_104(wire_con_in_stage2[104]), .outData_105(wire_con_in_stage2[105]), .outData_106(wire_con_in_stage2[106]), .outData_107(wire_con_in_stage2[107]), .outData_108(wire_con_in_stage2[108]), .outData_109(wire_con_in_stage2[109]), .outData_110(wire_con_in_stage2[110]), .outData_111(wire_con_in_stage2[111]), .outData_112(wire_con_in_stage2[112]), .outData_113(wire_con_in_stage2[113]), .outData_114(wire_con_in_stage2[114]), .outData_115(wire_con_in_stage2[115]), .outData_116(wire_con_in_stage2[116]), .outData_117(wire_con_in_stage2[117]), .outData_118(wire_con_in_stage2[118]), .outData_119(wire_con_in_stage2[119]), .outData_120(wire_con_in_stage2[120]), .outData_121(wire_con_in_stage2[121]), .outData_122(wire_con_in_stage2[122]), .outData_123(wire_con_in_stage2[123]), .outData_124(wire_con_in_stage2[124]), .outData_125(wire_con_in_stage2[125]), .outData_126(wire_con_in_stage2[126]), .outData_127(wire_con_in_stage2[127]), .outData_128(wire_con_in_stage2[128]), .outData_129(wire_con_in_stage2[129]), .outData_130(wire_con_in_stage2[130]), .outData_131(wire_con_in_stage2[131]), .outData_132(wire_con_in_stage2[132]), .outData_133(wire_con_in_stage2[133]), .outData_134(wire_con_in_stage2[134]), .outData_135(wire_con_in_stage2[135]), .outData_136(wire_con_in_stage2[136]), .outData_137(wire_con_in_stage2[137]), .outData_138(wire_con_in_stage2[138]), .outData_139(wire_con_in_stage2[139]), .outData_140(wire_con_in_stage2[140]), .outData_141(wire_con_in_stage2[141]), .outData_142(wire_con_in_stage2[142]), .outData_143(wire_con_in_stage2[143]), .outData_144(wire_con_in_stage2[144]), .outData_145(wire_con_in_stage2[145]), .outData_146(wire_con_in_stage2[146]), .outData_147(wire_con_in_stage2[147]), .outData_148(wire_con_in_stage2[148]), .outData_149(wire_con_in_stage2[149]), .outData_150(wire_con_in_stage2[150]), .outData_151(wire_con_in_stage2[151]), .outData_152(wire_con_in_stage2[152]), .outData_153(wire_con_in_stage2[153]), .outData_154(wire_con_in_stage2[154]), .outData_155(wire_con_in_stage2[155]), .outData_156(wire_con_in_stage2[156]), .outData_157(wire_con_in_stage2[157]), .outData_158(wire_con_in_stage2[158]), .outData_159(wire_con_in_stage2[159]), .outData_160(wire_con_in_stage2[160]), .outData_161(wire_con_in_stage2[161]), .outData_162(wire_con_in_stage2[162]), .outData_163(wire_con_in_stage2[163]), .outData_164(wire_con_in_stage2[164]), .outData_165(wire_con_in_stage2[165]), .outData_166(wire_con_in_stage2[166]), .outData_167(wire_con_in_stage2[167]), .outData_168(wire_con_in_stage2[168]), .outData_169(wire_con_in_stage2[169]), .outData_170(wire_con_in_stage2[170]), .outData_171(wire_con_in_stage2[171]), .outData_172(wire_con_in_stage2[172]), .outData_173(wire_con_in_stage2[173]), .outData_174(wire_con_in_stage2[174]), .outData_175(wire_con_in_stage2[175]), .outData_176(wire_con_in_stage2[176]), .outData_177(wire_con_in_stage2[177]), .outData_178(wire_con_in_stage2[178]), .outData_179(wire_con_in_stage2[179]), .outData_180(wire_con_in_stage2[180]), .outData_181(wire_con_in_stage2[181]), .outData_182(wire_con_in_stage2[182]), .outData_183(wire_con_in_stage2[183]), .outData_184(wire_con_in_stage2[184]), .outData_185(wire_con_in_stage2[185]), .outData_186(wire_con_in_stage2[186]), .outData_187(wire_con_in_stage2[187]), .outData_188(wire_con_in_stage2[188]), .outData_189(wire_con_in_stage2[189]), .outData_190(wire_con_in_stage2[190]), .outData_191(wire_con_in_stage2[191]), .outData_192(wire_con_in_stage2[192]), .outData_193(wire_con_in_stage2[193]), .outData_194(wire_con_in_stage2[194]), .outData_195(wire_con_in_stage2[195]), .outData_196(wire_con_in_stage2[196]), .outData_197(wire_con_in_stage2[197]), .outData_198(wire_con_in_stage2[198]), .outData_199(wire_con_in_stage2[199]), .outData_200(wire_con_in_stage2[200]), .outData_201(wire_con_in_stage2[201]), .outData_202(wire_con_in_stage2[202]), .outData_203(wire_con_in_stage2[203]), .outData_204(wire_con_in_stage2[204]), .outData_205(wire_con_in_stage2[205]), .outData_206(wire_con_in_stage2[206]), .outData_207(wire_con_in_stage2[207]), .outData_208(wire_con_in_stage2[208]), .outData_209(wire_con_in_stage2[209]), .outData_210(wire_con_in_stage2[210]), .outData_211(wire_con_in_stage2[211]), .outData_212(wire_con_in_stage2[212]), .outData_213(wire_con_in_stage2[213]), .outData_214(wire_con_in_stage2[214]), .outData_215(wire_con_in_stage2[215]), .outData_216(wire_con_in_stage2[216]), .outData_217(wire_con_in_stage2[217]), .outData_218(wire_con_in_stage2[218]), .outData_219(wire_con_in_stage2[219]), .outData_220(wire_con_in_stage2[220]), .outData_221(wire_con_in_stage2[221]), .outData_222(wire_con_in_stage2[222]), .outData_223(wire_con_in_stage2[223]), .outData_224(wire_con_in_stage2[224]), .outData_225(wire_con_in_stage2[225]), .outData_226(wire_con_in_stage2[226]), .outData_227(wire_con_in_stage2[227]), .outData_228(wire_con_in_stage2[228]), .outData_229(wire_con_in_stage2[229]), .outData_230(wire_con_in_stage2[230]), .outData_231(wire_con_in_stage2[231]), .outData_232(wire_con_in_stage2[232]), .outData_233(wire_con_in_stage2[233]), .outData_234(wire_con_in_stage2[234]), .outData_235(wire_con_in_stage2[235]), .outData_236(wire_con_in_stage2[236]), .outData_237(wire_con_in_stage2[237]), .outData_238(wire_con_in_stage2[238]), .outData_239(wire_con_in_stage2[239]), .outData_240(wire_con_in_stage2[240]), .outData_241(wire_con_in_stage2[241]), .outData_242(wire_con_in_stage2[242]), .outData_243(wire_con_in_stage2[243]), .outData_244(wire_con_in_stage2[244]), .outData_245(wire_con_in_stage2[245]), .outData_246(wire_con_in_stage2[246]), .outData_247(wire_con_in_stage2[247]), .outData_248(wire_con_in_stage2[248]), .outData_249(wire_con_in_stage2[249]), .outData_250(wire_con_in_stage2[250]), .outData_251(wire_con_in_stage2[251]), .outData_252(wire_con_in_stage2[252]), .outData_253(wire_con_in_stage2[253]), .outData_254(wire_con_in_stage2[254]), .outData_255(wire_con_in_stage2[255]), 
        .in_start(in_start_stage2), .out_start(con_in_start_stage2), .ctrl(wire_ctrl_stage2), .clk(clk), .rst(rst));
  
  wireCon_dp256_st2_L wire_stage_2(
        .inData_0(wire_con_in_stage2[0]), .inData_1(wire_con_in_stage2[1]), .inData_2(wire_con_in_stage2[2]), .inData_3(wire_con_in_stage2[3]), .inData_4(wire_con_in_stage2[4]), .inData_5(wire_con_in_stage2[5]), .inData_6(wire_con_in_stage2[6]), .inData_7(wire_con_in_stage2[7]), .inData_8(wire_con_in_stage2[8]), .inData_9(wire_con_in_stage2[9]), .inData_10(wire_con_in_stage2[10]), .inData_11(wire_con_in_stage2[11]), .inData_12(wire_con_in_stage2[12]), .inData_13(wire_con_in_stage2[13]), .inData_14(wire_con_in_stage2[14]), .inData_15(wire_con_in_stage2[15]), .inData_16(wire_con_in_stage2[16]), .inData_17(wire_con_in_stage2[17]), .inData_18(wire_con_in_stage2[18]), .inData_19(wire_con_in_stage2[19]), .inData_20(wire_con_in_stage2[20]), .inData_21(wire_con_in_stage2[21]), .inData_22(wire_con_in_stage2[22]), .inData_23(wire_con_in_stage2[23]), .inData_24(wire_con_in_stage2[24]), .inData_25(wire_con_in_stage2[25]), .inData_26(wire_con_in_stage2[26]), .inData_27(wire_con_in_stage2[27]), .inData_28(wire_con_in_stage2[28]), .inData_29(wire_con_in_stage2[29]), .inData_30(wire_con_in_stage2[30]), .inData_31(wire_con_in_stage2[31]), .inData_32(wire_con_in_stage2[32]), .inData_33(wire_con_in_stage2[33]), .inData_34(wire_con_in_stage2[34]), .inData_35(wire_con_in_stage2[35]), .inData_36(wire_con_in_stage2[36]), .inData_37(wire_con_in_stage2[37]), .inData_38(wire_con_in_stage2[38]), .inData_39(wire_con_in_stage2[39]), .inData_40(wire_con_in_stage2[40]), .inData_41(wire_con_in_stage2[41]), .inData_42(wire_con_in_stage2[42]), .inData_43(wire_con_in_stage2[43]), .inData_44(wire_con_in_stage2[44]), .inData_45(wire_con_in_stage2[45]), .inData_46(wire_con_in_stage2[46]), .inData_47(wire_con_in_stage2[47]), .inData_48(wire_con_in_stage2[48]), .inData_49(wire_con_in_stage2[49]), .inData_50(wire_con_in_stage2[50]), .inData_51(wire_con_in_stage2[51]), .inData_52(wire_con_in_stage2[52]), .inData_53(wire_con_in_stage2[53]), .inData_54(wire_con_in_stage2[54]), .inData_55(wire_con_in_stage2[55]), .inData_56(wire_con_in_stage2[56]), .inData_57(wire_con_in_stage2[57]), .inData_58(wire_con_in_stage2[58]), .inData_59(wire_con_in_stage2[59]), .inData_60(wire_con_in_stage2[60]), .inData_61(wire_con_in_stage2[61]), .inData_62(wire_con_in_stage2[62]), .inData_63(wire_con_in_stage2[63]), .inData_64(wire_con_in_stage2[64]), .inData_65(wire_con_in_stage2[65]), .inData_66(wire_con_in_stage2[66]), .inData_67(wire_con_in_stage2[67]), .inData_68(wire_con_in_stage2[68]), .inData_69(wire_con_in_stage2[69]), .inData_70(wire_con_in_stage2[70]), .inData_71(wire_con_in_stage2[71]), .inData_72(wire_con_in_stage2[72]), .inData_73(wire_con_in_stage2[73]), .inData_74(wire_con_in_stage2[74]), .inData_75(wire_con_in_stage2[75]), .inData_76(wire_con_in_stage2[76]), .inData_77(wire_con_in_stage2[77]), .inData_78(wire_con_in_stage2[78]), .inData_79(wire_con_in_stage2[79]), .inData_80(wire_con_in_stage2[80]), .inData_81(wire_con_in_stage2[81]), .inData_82(wire_con_in_stage2[82]), .inData_83(wire_con_in_stage2[83]), .inData_84(wire_con_in_stage2[84]), .inData_85(wire_con_in_stage2[85]), .inData_86(wire_con_in_stage2[86]), .inData_87(wire_con_in_stage2[87]), .inData_88(wire_con_in_stage2[88]), .inData_89(wire_con_in_stage2[89]), .inData_90(wire_con_in_stage2[90]), .inData_91(wire_con_in_stage2[91]), .inData_92(wire_con_in_stage2[92]), .inData_93(wire_con_in_stage2[93]), .inData_94(wire_con_in_stage2[94]), .inData_95(wire_con_in_stage2[95]), .inData_96(wire_con_in_stage2[96]), .inData_97(wire_con_in_stage2[97]), .inData_98(wire_con_in_stage2[98]), .inData_99(wire_con_in_stage2[99]), .inData_100(wire_con_in_stage2[100]), .inData_101(wire_con_in_stage2[101]), .inData_102(wire_con_in_stage2[102]), .inData_103(wire_con_in_stage2[103]), .inData_104(wire_con_in_stage2[104]), .inData_105(wire_con_in_stage2[105]), .inData_106(wire_con_in_stage2[106]), .inData_107(wire_con_in_stage2[107]), .inData_108(wire_con_in_stage2[108]), .inData_109(wire_con_in_stage2[109]), .inData_110(wire_con_in_stage2[110]), .inData_111(wire_con_in_stage2[111]), .inData_112(wire_con_in_stage2[112]), .inData_113(wire_con_in_stage2[113]), .inData_114(wire_con_in_stage2[114]), .inData_115(wire_con_in_stage2[115]), .inData_116(wire_con_in_stage2[116]), .inData_117(wire_con_in_stage2[117]), .inData_118(wire_con_in_stage2[118]), .inData_119(wire_con_in_stage2[119]), .inData_120(wire_con_in_stage2[120]), .inData_121(wire_con_in_stage2[121]), .inData_122(wire_con_in_stage2[122]), .inData_123(wire_con_in_stage2[123]), .inData_124(wire_con_in_stage2[124]), .inData_125(wire_con_in_stage2[125]), .inData_126(wire_con_in_stage2[126]), .inData_127(wire_con_in_stage2[127]), .inData_128(wire_con_in_stage2[128]), .inData_129(wire_con_in_stage2[129]), .inData_130(wire_con_in_stage2[130]), .inData_131(wire_con_in_stage2[131]), .inData_132(wire_con_in_stage2[132]), .inData_133(wire_con_in_stage2[133]), .inData_134(wire_con_in_stage2[134]), .inData_135(wire_con_in_stage2[135]), .inData_136(wire_con_in_stage2[136]), .inData_137(wire_con_in_stage2[137]), .inData_138(wire_con_in_stage2[138]), .inData_139(wire_con_in_stage2[139]), .inData_140(wire_con_in_stage2[140]), .inData_141(wire_con_in_stage2[141]), .inData_142(wire_con_in_stage2[142]), .inData_143(wire_con_in_stage2[143]), .inData_144(wire_con_in_stage2[144]), .inData_145(wire_con_in_stage2[145]), .inData_146(wire_con_in_stage2[146]), .inData_147(wire_con_in_stage2[147]), .inData_148(wire_con_in_stage2[148]), .inData_149(wire_con_in_stage2[149]), .inData_150(wire_con_in_stage2[150]), .inData_151(wire_con_in_stage2[151]), .inData_152(wire_con_in_stage2[152]), .inData_153(wire_con_in_stage2[153]), .inData_154(wire_con_in_stage2[154]), .inData_155(wire_con_in_stage2[155]), .inData_156(wire_con_in_stage2[156]), .inData_157(wire_con_in_stage2[157]), .inData_158(wire_con_in_stage2[158]), .inData_159(wire_con_in_stage2[159]), .inData_160(wire_con_in_stage2[160]), .inData_161(wire_con_in_stage2[161]), .inData_162(wire_con_in_stage2[162]), .inData_163(wire_con_in_stage2[163]), .inData_164(wire_con_in_stage2[164]), .inData_165(wire_con_in_stage2[165]), .inData_166(wire_con_in_stage2[166]), .inData_167(wire_con_in_stage2[167]), .inData_168(wire_con_in_stage2[168]), .inData_169(wire_con_in_stage2[169]), .inData_170(wire_con_in_stage2[170]), .inData_171(wire_con_in_stage2[171]), .inData_172(wire_con_in_stage2[172]), .inData_173(wire_con_in_stage2[173]), .inData_174(wire_con_in_stage2[174]), .inData_175(wire_con_in_stage2[175]), .inData_176(wire_con_in_stage2[176]), .inData_177(wire_con_in_stage2[177]), .inData_178(wire_con_in_stage2[178]), .inData_179(wire_con_in_stage2[179]), .inData_180(wire_con_in_stage2[180]), .inData_181(wire_con_in_stage2[181]), .inData_182(wire_con_in_stage2[182]), .inData_183(wire_con_in_stage2[183]), .inData_184(wire_con_in_stage2[184]), .inData_185(wire_con_in_stage2[185]), .inData_186(wire_con_in_stage2[186]), .inData_187(wire_con_in_stage2[187]), .inData_188(wire_con_in_stage2[188]), .inData_189(wire_con_in_stage2[189]), .inData_190(wire_con_in_stage2[190]), .inData_191(wire_con_in_stage2[191]), .inData_192(wire_con_in_stage2[192]), .inData_193(wire_con_in_stage2[193]), .inData_194(wire_con_in_stage2[194]), .inData_195(wire_con_in_stage2[195]), .inData_196(wire_con_in_stage2[196]), .inData_197(wire_con_in_stage2[197]), .inData_198(wire_con_in_stage2[198]), .inData_199(wire_con_in_stage2[199]), .inData_200(wire_con_in_stage2[200]), .inData_201(wire_con_in_stage2[201]), .inData_202(wire_con_in_stage2[202]), .inData_203(wire_con_in_stage2[203]), .inData_204(wire_con_in_stage2[204]), .inData_205(wire_con_in_stage2[205]), .inData_206(wire_con_in_stage2[206]), .inData_207(wire_con_in_stage2[207]), .inData_208(wire_con_in_stage2[208]), .inData_209(wire_con_in_stage2[209]), .inData_210(wire_con_in_stage2[210]), .inData_211(wire_con_in_stage2[211]), .inData_212(wire_con_in_stage2[212]), .inData_213(wire_con_in_stage2[213]), .inData_214(wire_con_in_stage2[214]), .inData_215(wire_con_in_stage2[215]), .inData_216(wire_con_in_stage2[216]), .inData_217(wire_con_in_stage2[217]), .inData_218(wire_con_in_stage2[218]), .inData_219(wire_con_in_stage2[219]), .inData_220(wire_con_in_stage2[220]), .inData_221(wire_con_in_stage2[221]), .inData_222(wire_con_in_stage2[222]), .inData_223(wire_con_in_stage2[223]), .inData_224(wire_con_in_stage2[224]), .inData_225(wire_con_in_stage2[225]), .inData_226(wire_con_in_stage2[226]), .inData_227(wire_con_in_stage2[227]), .inData_228(wire_con_in_stage2[228]), .inData_229(wire_con_in_stage2[229]), .inData_230(wire_con_in_stage2[230]), .inData_231(wire_con_in_stage2[231]), .inData_232(wire_con_in_stage2[232]), .inData_233(wire_con_in_stage2[233]), .inData_234(wire_con_in_stage2[234]), .inData_235(wire_con_in_stage2[235]), .inData_236(wire_con_in_stage2[236]), .inData_237(wire_con_in_stage2[237]), .inData_238(wire_con_in_stage2[238]), .inData_239(wire_con_in_stage2[239]), .inData_240(wire_con_in_stage2[240]), .inData_241(wire_con_in_stage2[241]), .inData_242(wire_con_in_stage2[242]), .inData_243(wire_con_in_stage2[243]), .inData_244(wire_con_in_stage2[244]), .inData_245(wire_con_in_stage2[245]), .inData_246(wire_con_in_stage2[246]), .inData_247(wire_con_in_stage2[247]), .inData_248(wire_con_in_stage2[248]), .inData_249(wire_con_in_stage2[249]), .inData_250(wire_con_in_stage2[250]), .inData_251(wire_con_in_stage2[251]), .inData_252(wire_con_in_stage2[252]), .inData_253(wire_con_in_stage2[253]), .inData_254(wire_con_in_stage2[254]), .inData_255(wire_con_in_stage2[255]), 
        .outData_0(wire_con_out_stage2[0]), .outData_1(wire_con_out_stage2[1]), .outData_2(wire_con_out_stage2[2]), .outData_3(wire_con_out_stage2[3]), .outData_4(wire_con_out_stage2[4]), .outData_5(wire_con_out_stage2[5]), .outData_6(wire_con_out_stage2[6]), .outData_7(wire_con_out_stage2[7]), .outData_8(wire_con_out_stage2[8]), .outData_9(wire_con_out_stage2[9]), .outData_10(wire_con_out_stage2[10]), .outData_11(wire_con_out_stage2[11]), .outData_12(wire_con_out_stage2[12]), .outData_13(wire_con_out_stage2[13]), .outData_14(wire_con_out_stage2[14]), .outData_15(wire_con_out_stage2[15]), .outData_16(wire_con_out_stage2[16]), .outData_17(wire_con_out_stage2[17]), .outData_18(wire_con_out_stage2[18]), .outData_19(wire_con_out_stage2[19]), .outData_20(wire_con_out_stage2[20]), .outData_21(wire_con_out_stage2[21]), .outData_22(wire_con_out_stage2[22]), .outData_23(wire_con_out_stage2[23]), .outData_24(wire_con_out_stage2[24]), .outData_25(wire_con_out_stage2[25]), .outData_26(wire_con_out_stage2[26]), .outData_27(wire_con_out_stage2[27]), .outData_28(wire_con_out_stage2[28]), .outData_29(wire_con_out_stage2[29]), .outData_30(wire_con_out_stage2[30]), .outData_31(wire_con_out_stage2[31]), .outData_32(wire_con_out_stage2[32]), .outData_33(wire_con_out_stage2[33]), .outData_34(wire_con_out_stage2[34]), .outData_35(wire_con_out_stage2[35]), .outData_36(wire_con_out_stage2[36]), .outData_37(wire_con_out_stage2[37]), .outData_38(wire_con_out_stage2[38]), .outData_39(wire_con_out_stage2[39]), .outData_40(wire_con_out_stage2[40]), .outData_41(wire_con_out_stage2[41]), .outData_42(wire_con_out_stage2[42]), .outData_43(wire_con_out_stage2[43]), .outData_44(wire_con_out_stage2[44]), .outData_45(wire_con_out_stage2[45]), .outData_46(wire_con_out_stage2[46]), .outData_47(wire_con_out_stage2[47]), .outData_48(wire_con_out_stage2[48]), .outData_49(wire_con_out_stage2[49]), .outData_50(wire_con_out_stage2[50]), .outData_51(wire_con_out_stage2[51]), .outData_52(wire_con_out_stage2[52]), .outData_53(wire_con_out_stage2[53]), .outData_54(wire_con_out_stage2[54]), .outData_55(wire_con_out_stage2[55]), .outData_56(wire_con_out_stage2[56]), .outData_57(wire_con_out_stage2[57]), .outData_58(wire_con_out_stage2[58]), .outData_59(wire_con_out_stage2[59]), .outData_60(wire_con_out_stage2[60]), .outData_61(wire_con_out_stage2[61]), .outData_62(wire_con_out_stage2[62]), .outData_63(wire_con_out_stage2[63]), .outData_64(wire_con_out_stage2[64]), .outData_65(wire_con_out_stage2[65]), .outData_66(wire_con_out_stage2[66]), .outData_67(wire_con_out_stage2[67]), .outData_68(wire_con_out_stage2[68]), .outData_69(wire_con_out_stage2[69]), .outData_70(wire_con_out_stage2[70]), .outData_71(wire_con_out_stage2[71]), .outData_72(wire_con_out_stage2[72]), .outData_73(wire_con_out_stage2[73]), .outData_74(wire_con_out_stage2[74]), .outData_75(wire_con_out_stage2[75]), .outData_76(wire_con_out_stage2[76]), .outData_77(wire_con_out_stage2[77]), .outData_78(wire_con_out_stage2[78]), .outData_79(wire_con_out_stage2[79]), .outData_80(wire_con_out_stage2[80]), .outData_81(wire_con_out_stage2[81]), .outData_82(wire_con_out_stage2[82]), .outData_83(wire_con_out_stage2[83]), .outData_84(wire_con_out_stage2[84]), .outData_85(wire_con_out_stage2[85]), .outData_86(wire_con_out_stage2[86]), .outData_87(wire_con_out_stage2[87]), .outData_88(wire_con_out_stage2[88]), .outData_89(wire_con_out_stage2[89]), .outData_90(wire_con_out_stage2[90]), .outData_91(wire_con_out_stage2[91]), .outData_92(wire_con_out_stage2[92]), .outData_93(wire_con_out_stage2[93]), .outData_94(wire_con_out_stage2[94]), .outData_95(wire_con_out_stage2[95]), .outData_96(wire_con_out_stage2[96]), .outData_97(wire_con_out_stage2[97]), .outData_98(wire_con_out_stage2[98]), .outData_99(wire_con_out_stage2[99]), .outData_100(wire_con_out_stage2[100]), .outData_101(wire_con_out_stage2[101]), .outData_102(wire_con_out_stage2[102]), .outData_103(wire_con_out_stage2[103]), .outData_104(wire_con_out_stage2[104]), .outData_105(wire_con_out_stage2[105]), .outData_106(wire_con_out_stage2[106]), .outData_107(wire_con_out_stage2[107]), .outData_108(wire_con_out_stage2[108]), .outData_109(wire_con_out_stage2[109]), .outData_110(wire_con_out_stage2[110]), .outData_111(wire_con_out_stage2[111]), .outData_112(wire_con_out_stage2[112]), .outData_113(wire_con_out_stage2[113]), .outData_114(wire_con_out_stage2[114]), .outData_115(wire_con_out_stage2[115]), .outData_116(wire_con_out_stage2[116]), .outData_117(wire_con_out_stage2[117]), .outData_118(wire_con_out_stage2[118]), .outData_119(wire_con_out_stage2[119]), .outData_120(wire_con_out_stage2[120]), .outData_121(wire_con_out_stage2[121]), .outData_122(wire_con_out_stage2[122]), .outData_123(wire_con_out_stage2[123]), .outData_124(wire_con_out_stage2[124]), .outData_125(wire_con_out_stage2[125]), .outData_126(wire_con_out_stage2[126]), .outData_127(wire_con_out_stage2[127]), .outData_128(wire_con_out_stage2[128]), .outData_129(wire_con_out_stage2[129]), .outData_130(wire_con_out_stage2[130]), .outData_131(wire_con_out_stage2[131]), .outData_132(wire_con_out_stage2[132]), .outData_133(wire_con_out_stage2[133]), .outData_134(wire_con_out_stage2[134]), .outData_135(wire_con_out_stage2[135]), .outData_136(wire_con_out_stage2[136]), .outData_137(wire_con_out_stage2[137]), .outData_138(wire_con_out_stage2[138]), .outData_139(wire_con_out_stage2[139]), .outData_140(wire_con_out_stage2[140]), .outData_141(wire_con_out_stage2[141]), .outData_142(wire_con_out_stage2[142]), .outData_143(wire_con_out_stage2[143]), .outData_144(wire_con_out_stage2[144]), .outData_145(wire_con_out_stage2[145]), .outData_146(wire_con_out_stage2[146]), .outData_147(wire_con_out_stage2[147]), .outData_148(wire_con_out_stage2[148]), .outData_149(wire_con_out_stage2[149]), .outData_150(wire_con_out_stage2[150]), .outData_151(wire_con_out_stage2[151]), .outData_152(wire_con_out_stage2[152]), .outData_153(wire_con_out_stage2[153]), .outData_154(wire_con_out_stage2[154]), .outData_155(wire_con_out_stage2[155]), .outData_156(wire_con_out_stage2[156]), .outData_157(wire_con_out_stage2[157]), .outData_158(wire_con_out_stage2[158]), .outData_159(wire_con_out_stage2[159]), .outData_160(wire_con_out_stage2[160]), .outData_161(wire_con_out_stage2[161]), .outData_162(wire_con_out_stage2[162]), .outData_163(wire_con_out_stage2[163]), .outData_164(wire_con_out_stage2[164]), .outData_165(wire_con_out_stage2[165]), .outData_166(wire_con_out_stage2[166]), .outData_167(wire_con_out_stage2[167]), .outData_168(wire_con_out_stage2[168]), .outData_169(wire_con_out_stage2[169]), .outData_170(wire_con_out_stage2[170]), .outData_171(wire_con_out_stage2[171]), .outData_172(wire_con_out_stage2[172]), .outData_173(wire_con_out_stage2[173]), .outData_174(wire_con_out_stage2[174]), .outData_175(wire_con_out_stage2[175]), .outData_176(wire_con_out_stage2[176]), .outData_177(wire_con_out_stage2[177]), .outData_178(wire_con_out_stage2[178]), .outData_179(wire_con_out_stage2[179]), .outData_180(wire_con_out_stage2[180]), .outData_181(wire_con_out_stage2[181]), .outData_182(wire_con_out_stage2[182]), .outData_183(wire_con_out_stage2[183]), .outData_184(wire_con_out_stage2[184]), .outData_185(wire_con_out_stage2[185]), .outData_186(wire_con_out_stage2[186]), .outData_187(wire_con_out_stage2[187]), .outData_188(wire_con_out_stage2[188]), .outData_189(wire_con_out_stage2[189]), .outData_190(wire_con_out_stage2[190]), .outData_191(wire_con_out_stage2[191]), .outData_192(wire_con_out_stage2[192]), .outData_193(wire_con_out_stage2[193]), .outData_194(wire_con_out_stage2[194]), .outData_195(wire_con_out_stage2[195]), .outData_196(wire_con_out_stage2[196]), .outData_197(wire_con_out_stage2[197]), .outData_198(wire_con_out_stage2[198]), .outData_199(wire_con_out_stage2[199]), .outData_200(wire_con_out_stage2[200]), .outData_201(wire_con_out_stage2[201]), .outData_202(wire_con_out_stage2[202]), .outData_203(wire_con_out_stage2[203]), .outData_204(wire_con_out_stage2[204]), .outData_205(wire_con_out_stage2[205]), .outData_206(wire_con_out_stage2[206]), .outData_207(wire_con_out_stage2[207]), .outData_208(wire_con_out_stage2[208]), .outData_209(wire_con_out_stage2[209]), .outData_210(wire_con_out_stage2[210]), .outData_211(wire_con_out_stage2[211]), .outData_212(wire_con_out_stage2[212]), .outData_213(wire_con_out_stage2[213]), .outData_214(wire_con_out_stage2[214]), .outData_215(wire_con_out_stage2[215]), .outData_216(wire_con_out_stage2[216]), .outData_217(wire_con_out_stage2[217]), .outData_218(wire_con_out_stage2[218]), .outData_219(wire_con_out_stage2[219]), .outData_220(wire_con_out_stage2[220]), .outData_221(wire_con_out_stage2[221]), .outData_222(wire_con_out_stage2[222]), .outData_223(wire_con_out_stage2[223]), .outData_224(wire_con_out_stage2[224]), .outData_225(wire_con_out_stage2[225]), .outData_226(wire_con_out_stage2[226]), .outData_227(wire_con_out_stage2[227]), .outData_228(wire_con_out_stage2[228]), .outData_229(wire_con_out_stage2[229]), .outData_230(wire_con_out_stage2[230]), .outData_231(wire_con_out_stage2[231]), .outData_232(wire_con_out_stage2[232]), .outData_233(wire_con_out_stage2[233]), .outData_234(wire_con_out_stage2[234]), .outData_235(wire_con_out_stage2[235]), .outData_236(wire_con_out_stage2[236]), .outData_237(wire_con_out_stage2[237]), .outData_238(wire_con_out_stage2[238]), .outData_239(wire_con_out_stage2[239]), .outData_240(wire_con_out_stage2[240]), .outData_241(wire_con_out_stage2[241]), .outData_242(wire_con_out_stage2[242]), .outData_243(wire_con_out_stage2[243]), .outData_244(wire_con_out_stage2[244]), .outData_245(wire_con_out_stage2[245]), .outData_246(wire_con_out_stage2[246]), .outData_247(wire_con_out_stage2[247]), .outData_248(wire_con_out_stage2[248]), .outData_249(wire_con_out_stage2[249]), .outData_250(wire_con_out_stage2[250]), .outData_251(wire_con_out_stage2[251]), .outData_252(wire_con_out_stage2[252]), .outData_253(wire_con_out_stage2[253]), .outData_254(wire_con_out_stage2[254]), .outData_255(wire_con_out_stage2[255]), 
        .in_start(con_in_start_stage2), .out_start(in_start_stage3), .clk(clk), .rst(rst)); 

  
  assign wire_ctrl_stage2[0] = counter_w[5]; 
  assign wire_ctrl_stage2[1] = counter_w[5]; 
  assign wire_ctrl_stage2[2] = counter_w[5]; 
  assign wire_ctrl_stage2[3] = counter_w[5]; 
  assign wire_ctrl_stage2[4] = counter_w[5]; 
  assign wire_ctrl_stage2[5] = counter_w[5]; 
  assign wire_ctrl_stage2[6] = counter_w[5]; 
  assign wire_ctrl_stage2[7] = counter_w[5]; 
  assign wire_ctrl_stage2[8] = counter_w[5]; 
  assign wire_ctrl_stage2[9] = counter_w[5]; 
  assign wire_ctrl_stage2[10] = counter_w[5]; 
  assign wire_ctrl_stage2[11] = counter_w[5]; 
  assign wire_ctrl_stage2[12] = counter_w[5]; 
  assign wire_ctrl_stage2[13] = counter_w[5]; 
  assign wire_ctrl_stage2[14] = counter_w[5]; 
  assign wire_ctrl_stage2[15] = counter_w[5]; 
  assign wire_ctrl_stage2[16] = counter_w[5]; 
  assign wire_ctrl_stage2[17] = counter_w[5]; 
  assign wire_ctrl_stage2[18] = counter_w[5]; 
  assign wire_ctrl_stage2[19] = counter_w[5]; 
  assign wire_ctrl_stage2[20] = counter_w[5]; 
  assign wire_ctrl_stage2[21] = counter_w[5]; 
  assign wire_ctrl_stage2[22] = counter_w[5]; 
  assign wire_ctrl_stage2[23] = counter_w[5]; 
  assign wire_ctrl_stage2[24] = counter_w[5]; 
  assign wire_ctrl_stage2[25] = counter_w[5]; 
  assign wire_ctrl_stage2[26] = counter_w[5]; 
  assign wire_ctrl_stage2[27] = counter_w[5]; 
  assign wire_ctrl_stage2[28] = counter_w[5]; 
  assign wire_ctrl_stage2[29] = counter_w[5]; 
  assign wire_ctrl_stage2[30] = counter_w[5]; 
  assign wire_ctrl_stage2[31] = counter_w[5]; 
  assign wire_ctrl_stage2[32] = counter_w[5]; 
  assign wire_ctrl_stage2[33] = counter_w[5]; 
  assign wire_ctrl_stage2[34] = counter_w[5]; 
  assign wire_ctrl_stage2[35] = counter_w[5]; 
  assign wire_ctrl_stage2[36] = counter_w[5]; 
  assign wire_ctrl_stage2[37] = counter_w[5]; 
  assign wire_ctrl_stage2[38] = counter_w[5]; 
  assign wire_ctrl_stage2[39] = counter_w[5]; 
  assign wire_ctrl_stage2[40] = counter_w[5]; 
  assign wire_ctrl_stage2[41] = counter_w[5]; 
  assign wire_ctrl_stage2[42] = counter_w[5]; 
  assign wire_ctrl_stage2[43] = counter_w[5]; 
  assign wire_ctrl_stage2[44] = counter_w[5]; 
  assign wire_ctrl_stage2[45] = counter_w[5]; 
  assign wire_ctrl_stage2[46] = counter_w[5]; 
  assign wire_ctrl_stage2[47] = counter_w[5]; 
  assign wire_ctrl_stage2[48] = counter_w[5]; 
  assign wire_ctrl_stage2[49] = counter_w[5]; 
  assign wire_ctrl_stage2[50] = counter_w[5]; 
  assign wire_ctrl_stage2[51] = counter_w[5]; 
  assign wire_ctrl_stage2[52] = counter_w[5]; 
  assign wire_ctrl_stage2[53] = counter_w[5]; 
  assign wire_ctrl_stage2[54] = counter_w[5]; 
  assign wire_ctrl_stage2[55] = counter_w[5]; 
  assign wire_ctrl_stage2[56] = counter_w[5]; 
  assign wire_ctrl_stage2[57] = counter_w[5]; 
  assign wire_ctrl_stage2[58] = counter_w[5]; 
  assign wire_ctrl_stage2[59] = counter_w[5]; 
  assign wire_ctrl_stage2[60] = counter_w[5]; 
  assign wire_ctrl_stage2[61] = counter_w[5]; 
  assign wire_ctrl_stage2[62] = counter_w[5]; 
  assign wire_ctrl_stage2[63] = counter_w[5]; 
  assign wire_ctrl_stage2[64] = counter_w[5]; 
  assign wire_ctrl_stage2[65] = counter_w[5]; 
  assign wire_ctrl_stage2[66] = counter_w[5]; 
  assign wire_ctrl_stage2[67] = counter_w[5]; 
  assign wire_ctrl_stage2[68] = counter_w[5]; 
  assign wire_ctrl_stage2[69] = counter_w[5]; 
  assign wire_ctrl_stage2[70] = counter_w[5]; 
  assign wire_ctrl_stage2[71] = counter_w[5]; 
  assign wire_ctrl_stage2[72] = counter_w[5]; 
  assign wire_ctrl_stage2[73] = counter_w[5]; 
  assign wire_ctrl_stage2[74] = counter_w[5]; 
  assign wire_ctrl_stage2[75] = counter_w[5]; 
  assign wire_ctrl_stage2[76] = counter_w[5]; 
  assign wire_ctrl_stage2[77] = counter_w[5]; 
  assign wire_ctrl_stage2[78] = counter_w[5]; 
  assign wire_ctrl_stage2[79] = counter_w[5]; 
  assign wire_ctrl_stage2[80] = counter_w[5]; 
  assign wire_ctrl_stage2[81] = counter_w[5]; 
  assign wire_ctrl_stage2[82] = counter_w[5]; 
  assign wire_ctrl_stage2[83] = counter_w[5]; 
  assign wire_ctrl_stage2[84] = counter_w[5]; 
  assign wire_ctrl_stage2[85] = counter_w[5]; 
  assign wire_ctrl_stage2[86] = counter_w[5]; 
  assign wire_ctrl_stage2[87] = counter_w[5]; 
  assign wire_ctrl_stage2[88] = counter_w[5]; 
  assign wire_ctrl_stage2[89] = counter_w[5]; 
  assign wire_ctrl_stage2[90] = counter_w[5]; 
  assign wire_ctrl_stage2[91] = counter_w[5]; 
  assign wire_ctrl_stage2[92] = counter_w[5]; 
  assign wire_ctrl_stage2[93] = counter_w[5]; 
  assign wire_ctrl_stage2[94] = counter_w[5]; 
  assign wire_ctrl_stage2[95] = counter_w[5]; 
  assign wire_ctrl_stage2[96] = counter_w[5]; 
  assign wire_ctrl_stage2[97] = counter_w[5]; 
  assign wire_ctrl_stage2[98] = counter_w[5]; 
  assign wire_ctrl_stage2[99] = counter_w[5]; 
  assign wire_ctrl_stage2[100] = counter_w[5]; 
  assign wire_ctrl_stage2[101] = counter_w[5]; 
  assign wire_ctrl_stage2[102] = counter_w[5]; 
  assign wire_ctrl_stage2[103] = counter_w[5]; 
  assign wire_ctrl_stage2[104] = counter_w[5]; 
  assign wire_ctrl_stage2[105] = counter_w[5]; 
  assign wire_ctrl_stage2[106] = counter_w[5]; 
  assign wire_ctrl_stage2[107] = counter_w[5]; 
  assign wire_ctrl_stage2[108] = counter_w[5]; 
  assign wire_ctrl_stage2[109] = counter_w[5]; 
  assign wire_ctrl_stage2[110] = counter_w[5]; 
  assign wire_ctrl_stage2[111] = counter_w[5]; 
  assign wire_ctrl_stage2[112] = counter_w[5]; 
  assign wire_ctrl_stage2[113] = counter_w[5]; 
  assign wire_ctrl_stage2[114] = counter_w[5]; 
  assign wire_ctrl_stage2[115] = counter_w[5]; 
  assign wire_ctrl_stage2[116] = counter_w[5]; 
  assign wire_ctrl_stage2[117] = counter_w[5]; 
  assign wire_ctrl_stage2[118] = counter_w[5]; 
  assign wire_ctrl_stage2[119] = counter_w[5]; 
  assign wire_ctrl_stage2[120] = counter_w[5]; 
  assign wire_ctrl_stage2[121] = counter_w[5]; 
  assign wire_ctrl_stage2[122] = counter_w[5]; 
  assign wire_ctrl_stage2[123] = counter_w[5]; 
  assign wire_ctrl_stage2[124] = counter_w[5]; 
  assign wire_ctrl_stage2[125] = counter_w[5]; 
  assign wire_ctrl_stage2[126] = counter_w[5]; 
  assign wire_ctrl_stage2[127] = counter_w[5]; 
  wire [DATA_WIDTH-1:0] wire_con_in_stage3[255:0];
  wire [DATA_WIDTH-1:0] wire_con_out_stage3[255:0];
  wire [127:0] wire_ctrl_stage3;

  switches_stage_st3_0_L switch_stage_3(
        .inData_0(wire_con_out_stage2[0]), .inData_1(wire_con_out_stage2[1]), .inData_2(wire_con_out_stage2[2]), .inData_3(wire_con_out_stage2[3]), .inData_4(wire_con_out_stage2[4]), .inData_5(wire_con_out_stage2[5]), .inData_6(wire_con_out_stage2[6]), .inData_7(wire_con_out_stage2[7]), .inData_8(wire_con_out_stage2[8]), .inData_9(wire_con_out_stage2[9]), .inData_10(wire_con_out_stage2[10]), .inData_11(wire_con_out_stage2[11]), .inData_12(wire_con_out_stage2[12]), .inData_13(wire_con_out_stage2[13]), .inData_14(wire_con_out_stage2[14]), .inData_15(wire_con_out_stage2[15]), .inData_16(wire_con_out_stage2[16]), .inData_17(wire_con_out_stage2[17]), .inData_18(wire_con_out_stage2[18]), .inData_19(wire_con_out_stage2[19]), .inData_20(wire_con_out_stage2[20]), .inData_21(wire_con_out_stage2[21]), .inData_22(wire_con_out_stage2[22]), .inData_23(wire_con_out_stage2[23]), .inData_24(wire_con_out_stage2[24]), .inData_25(wire_con_out_stage2[25]), .inData_26(wire_con_out_stage2[26]), .inData_27(wire_con_out_stage2[27]), .inData_28(wire_con_out_stage2[28]), .inData_29(wire_con_out_stage2[29]), .inData_30(wire_con_out_stage2[30]), .inData_31(wire_con_out_stage2[31]), .inData_32(wire_con_out_stage2[32]), .inData_33(wire_con_out_stage2[33]), .inData_34(wire_con_out_stage2[34]), .inData_35(wire_con_out_stage2[35]), .inData_36(wire_con_out_stage2[36]), .inData_37(wire_con_out_stage2[37]), .inData_38(wire_con_out_stage2[38]), .inData_39(wire_con_out_stage2[39]), .inData_40(wire_con_out_stage2[40]), .inData_41(wire_con_out_stage2[41]), .inData_42(wire_con_out_stage2[42]), .inData_43(wire_con_out_stage2[43]), .inData_44(wire_con_out_stage2[44]), .inData_45(wire_con_out_stage2[45]), .inData_46(wire_con_out_stage2[46]), .inData_47(wire_con_out_stage2[47]), .inData_48(wire_con_out_stage2[48]), .inData_49(wire_con_out_stage2[49]), .inData_50(wire_con_out_stage2[50]), .inData_51(wire_con_out_stage2[51]), .inData_52(wire_con_out_stage2[52]), .inData_53(wire_con_out_stage2[53]), .inData_54(wire_con_out_stage2[54]), .inData_55(wire_con_out_stage2[55]), .inData_56(wire_con_out_stage2[56]), .inData_57(wire_con_out_stage2[57]), .inData_58(wire_con_out_stage2[58]), .inData_59(wire_con_out_stage2[59]), .inData_60(wire_con_out_stage2[60]), .inData_61(wire_con_out_stage2[61]), .inData_62(wire_con_out_stage2[62]), .inData_63(wire_con_out_stage2[63]), .inData_64(wire_con_out_stage2[64]), .inData_65(wire_con_out_stage2[65]), .inData_66(wire_con_out_stage2[66]), .inData_67(wire_con_out_stage2[67]), .inData_68(wire_con_out_stage2[68]), .inData_69(wire_con_out_stage2[69]), .inData_70(wire_con_out_stage2[70]), .inData_71(wire_con_out_stage2[71]), .inData_72(wire_con_out_stage2[72]), .inData_73(wire_con_out_stage2[73]), .inData_74(wire_con_out_stage2[74]), .inData_75(wire_con_out_stage2[75]), .inData_76(wire_con_out_stage2[76]), .inData_77(wire_con_out_stage2[77]), .inData_78(wire_con_out_stage2[78]), .inData_79(wire_con_out_stage2[79]), .inData_80(wire_con_out_stage2[80]), .inData_81(wire_con_out_stage2[81]), .inData_82(wire_con_out_stage2[82]), .inData_83(wire_con_out_stage2[83]), .inData_84(wire_con_out_stage2[84]), .inData_85(wire_con_out_stage2[85]), .inData_86(wire_con_out_stage2[86]), .inData_87(wire_con_out_stage2[87]), .inData_88(wire_con_out_stage2[88]), .inData_89(wire_con_out_stage2[89]), .inData_90(wire_con_out_stage2[90]), .inData_91(wire_con_out_stage2[91]), .inData_92(wire_con_out_stage2[92]), .inData_93(wire_con_out_stage2[93]), .inData_94(wire_con_out_stage2[94]), .inData_95(wire_con_out_stage2[95]), .inData_96(wire_con_out_stage2[96]), .inData_97(wire_con_out_stage2[97]), .inData_98(wire_con_out_stage2[98]), .inData_99(wire_con_out_stage2[99]), .inData_100(wire_con_out_stage2[100]), .inData_101(wire_con_out_stage2[101]), .inData_102(wire_con_out_stage2[102]), .inData_103(wire_con_out_stage2[103]), .inData_104(wire_con_out_stage2[104]), .inData_105(wire_con_out_stage2[105]), .inData_106(wire_con_out_stage2[106]), .inData_107(wire_con_out_stage2[107]), .inData_108(wire_con_out_stage2[108]), .inData_109(wire_con_out_stage2[109]), .inData_110(wire_con_out_stage2[110]), .inData_111(wire_con_out_stage2[111]), .inData_112(wire_con_out_stage2[112]), .inData_113(wire_con_out_stage2[113]), .inData_114(wire_con_out_stage2[114]), .inData_115(wire_con_out_stage2[115]), .inData_116(wire_con_out_stage2[116]), .inData_117(wire_con_out_stage2[117]), .inData_118(wire_con_out_stage2[118]), .inData_119(wire_con_out_stage2[119]), .inData_120(wire_con_out_stage2[120]), .inData_121(wire_con_out_stage2[121]), .inData_122(wire_con_out_stage2[122]), .inData_123(wire_con_out_stage2[123]), .inData_124(wire_con_out_stage2[124]), .inData_125(wire_con_out_stage2[125]), .inData_126(wire_con_out_stage2[126]), .inData_127(wire_con_out_stage2[127]), .inData_128(wire_con_out_stage2[128]), .inData_129(wire_con_out_stage2[129]), .inData_130(wire_con_out_stage2[130]), .inData_131(wire_con_out_stage2[131]), .inData_132(wire_con_out_stage2[132]), .inData_133(wire_con_out_stage2[133]), .inData_134(wire_con_out_stage2[134]), .inData_135(wire_con_out_stage2[135]), .inData_136(wire_con_out_stage2[136]), .inData_137(wire_con_out_stage2[137]), .inData_138(wire_con_out_stage2[138]), .inData_139(wire_con_out_stage2[139]), .inData_140(wire_con_out_stage2[140]), .inData_141(wire_con_out_stage2[141]), .inData_142(wire_con_out_stage2[142]), .inData_143(wire_con_out_stage2[143]), .inData_144(wire_con_out_stage2[144]), .inData_145(wire_con_out_stage2[145]), .inData_146(wire_con_out_stage2[146]), .inData_147(wire_con_out_stage2[147]), .inData_148(wire_con_out_stage2[148]), .inData_149(wire_con_out_stage2[149]), .inData_150(wire_con_out_stage2[150]), .inData_151(wire_con_out_stage2[151]), .inData_152(wire_con_out_stage2[152]), .inData_153(wire_con_out_stage2[153]), .inData_154(wire_con_out_stage2[154]), .inData_155(wire_con_out_stage2[155]), .inData_156(wire_con_out_stage2[156]), .inData_157(wire_con_out_stage2[157]), .inData_158(wire_con_out_stage2[158]), .inData_159(wire_con_out_stage2[159]), .inData_160(wire_con_out_stage2[160]), .inData_161(wire_con_out_stage2[161]), .inData_162(wire_con_out_stage2[162]), .inData_163(wire_con_out_stage2[163]), .inData_164(wire_con_out_stage2[164]), .inData_165(wire_con_out_stage2[165]), .inData_166(wire_con_out_stage2[166]), .inData_167(wire_con_out_stage2[167]), .inData_168(wire_con_out_stage2[168]), .inData_169(wire_con_out_stage2[169]), .inData_170(wire_con_out_stage2[170]), .inData_171(wire_con_out_stage2[171]), .inData_172(wire_con_out_stage2[172]), .inData_173(wire_con_out_stage2[173]), .inData_174(wire_con_out_stage2[174]), .inData_175(wire_con_out_stage2[175]), .inData_176(wire_con_out_stage2[176]), .inData_177(wire_con_out_stage2[177]), .inData_178(wire_con_out_stage2[178]), .inData_179(wire_con_out_stage2[179]), .inData_180(wire_con_out_stage2[180]), .inData_181(wire_con_out_stage2[181]), .inData_182(wire_con_out_stage2[182]), .inData_183(wire_con_out_stage2[183]), .inData_184(wire_con_out_stage2[184]), .inData_185(wire_con_out_stage2[185]), .inData_186(wire_con_out_stage2[186]), .inData_187(wire_con_out_stage2[187]), .inData_188(wire_con_out_stage2[188]), .inData_189(wire_con_out_stage2[189]), .inData_190(wire_con_out_stage2[190]), .inData_191(wire_con_out_stage2[191]), .inData_192(wire_con_out_stage2[192]), .inData_193(wire_con_out_stage2[193]), .inData_194(wire_con_out_stage2[194]), .inData_195(wire_con_out_stage2[195]), .inData_196(wire_con_out_stage2[196]), .inData_197(wire_con_out_stage2[197]), .inData_198(wire_con_out_stage2[198]), .inData_199(wire_con_out_stage2[199]), .inData_200(wire_con_out_stage2[200]), .inData_201(wire_con_out_stage2[201]), .inData_202(wire_con_out_stage2[202]), .inData_203(wire_con_out_stage2[203]), .inData_204(wire_con_out_stage2[204]), .inData_205(wire_con_out_stage2[205]), .inData_206(wire_con_out_stage2[206]), .inData_207(wire_con_out_stage2[207]), .inData_208(wire_con_out_stage2[208]), .inData_209(wire_con_out_stage2[209]), .inData_210(wire_con_out_stage2[210]), .inData_211(wire_con_out_stage2[211]), .inData_212(wire_con_out_stage2[212]), .inData_213(wire_con_out_stage2[213]), .inData_214(wire_con_out_stage2[214]), .inData_215(wire_con_out_stage2[215]), .inData_216(wire_con_out_stage2[216]), .inData_217(wire_con_out_stage2[217]), .inData_218(wire_con_out_stage2[218]), .inData_219(wire_con_out_stage2[219]), .inData_220(wire_con_out_stage2[220]), .inData_221(wire_con_out_stage2[221]), .inData_222(wire_con_out_stage2[222]), .inData_223(wire_con_out_stage2[223]), .inData_224(wire_con_out_stage2[224]), .inData_225(wire_con_out_stage2[225]), .inData_226(wire_con_out_stage2[226]), .inData_227(wire_con_out_stage2[227]), .inData_228(wire_con_out_stage2[228]), .inData_229(wire_con_out_stage2[229]), .inData_230(wire_con_out_stage2[230]), .inData_231(wire_con_out_stage2[231]), .inData_232(wire_con_out_stage2[232]), .inData_233(wire_con_out_stage2[233]), .inData_234(wire_con_out_stage2[234]), .inData_235(wire_con_out_stage2[235]), .inData_236(wire_con_out_stage2[236]), .inData_237(wire_con_out_stage2[237]), .inData_238(wire_con_out_stage2[238]), .inData_239(wire_con_out_stage2[239]), .inData_240(wire_con_out_stage2[240]), .inData_241(wire_con_out_stage2[241]), .inData_242(wire_con_out_stage2[242]), .inData_243(wire_con_out_stage2[243]), .inData_244(wire_con_out_stage2[244]), .inData_245(wire_con_out_stage2[245]), .inData_246(wire_con_out_stage2[246]), .inData_247(wire_con_out_stage2[247]), .inData_248(wire_con_out_stage2[248]), .inData_249(wire_con_out_stage2[249]), .inData_250(wire_con_out_stage2[250]), .inData_251(wire_con_out_stage2[251]), .inData_252(wire_con_out_stage2[252]), .inData_253(wire_con_out_stage2[253]), .inData_254(wire_con_out_stage2[254]), .inData_255(wire_con_out_stage2[255]), 
        .outData_0(wire_con_in_stage3[0]), .outData_1(wire_con_in_stage3[1]), .outData_2(wire_con_in_stage3[2]), .outData_3(wire_con_in_stage3[3]), .outData_4(wire_con_in_stage3[4]), .outData_5(wire_con_in_stage3[5]), .outData_6(wire_con_in_stage3[6]), .outData_7(wire_con_in_stage3[7]), .outData_8(wire_con_in_stage3[8]), .outData_9(wire_con_in_stage3[9]), .outData_10(wire_con_in_stage3[10]), .outData_11(wire_con_in_stage3[11]), .outData_12(wire_con_in_stage3[12]), .outData_13(wire_con_in_stage3[13]), .outData_14(wire_con_in_stage3[14]), .outData_15(wire_con_in_stage3[15]), .outData_16(wire_con_in_stage3[16]), .outData_17(wire_con_in_stage3[17]), .outData_18(wire_con_in_stage3[18]), .outData_19(wire_con_in_stage3[19]), .outData_20(wire_con_in_stage3[20]), .outData_21(wire_con_in_stage3[21]), .outData_22(wire_con_in_stage3[22]), .outData_23(wire_con_in_stage3[23]), .outData_24(wire_con_in_stage3[24]), .outData_25(wire_con_in_stage3[25]), .outData_26(wire_con_in_stage3[26]), .outData_27(wire_con_in_stage3[27]), .outData_28(wire_con_in_stage3[28]), .outData_29(wire_con_in_stage3[29]), .outData_30(wire_con_in_stage3[30]), .outData_31(wire_con_in_stage3[31]), .outData_32(wire_con_in_stage3[32]), .outData_33(wire_con_in_stage3[33]), .outData_34(wire_con_in_stage3[34]), .outData_35(wire_con_in_stage3[35]), .outData_36(wire_con_in_stage3[36]), .outData_37(wire_con_in_stage3[37]), .outData_38(wire_con_in_stage3[38]), .outData_39(wire_con_in_stage3[39]), .outData_40(wire_con_in_stage3[40]), .outData_41(wire_con_in_stage3[41]), .outData_42(wire_con_in_stage3[42]), .outData_43(wire_con_in_stage3[43]), .outData_44(wire_con_in_stage3[44]), .outData_45(wire_con_in_stage3[45]), .outData_46(wire_con_in_stage3[46]), .outData_47(wire_con_in_stage3[47]), .outData_48(wire_con_in_stage3[48]), .outData_49(wire_con_in_stage3[49]), .outData_50(wire_con_in_stage3[50]), .outData_51(wire_con_in_stage3[51]), .outData_52(wire_con_in_stage3[52]), .outData_53(wire_con_in_stage3[53]), .outData_54(wire_con_in_stage3[54]), .outData_55(wire_con_in_stage3[55]), .outData_56(wire_con_in_stage3[56]), .outData_57(wire_con_in_stage3[57]), .outData_58(wire_con_in_stage3[58]), .outData_59(wire_con_in_stage3[59]), .outData_60(wire_con_in_stage3[60]), .outData_61(wire_con_in_stage3[61]), .outData_62(wire_con_in_stage3[62]), .outData_63(wire_con_in_stage3[63]), .outData_64(wire_con_in_stage3[64]), .outData_65(wire_con_in_stage3[65]), .outData_66(wire_con_in_stage3[66]), .outData_67(wire_con_in_stage3[67]), .outData_68(wire_con_in_stage3[68]), .outData_69(wire_con_in_stage3[69]), .outData_70(wire_con_in_stage3[70]), .outData_71(wire_con_in_stage3[71]), .outData_72(wire_con_in_stage3[72]), .outData_73(wire_con_in_stage3[73]), .outData_74(wire_con_in_stage3[74]), .outData_75(wire_con_in_stage3[75]), .outData_76(wire_con_in_stage3[76]), .outData_77(wire_con_in_stage3[77]), .outData_78(wire_con_in_stage3[78]), .outData_79(wire_con_in_stage3[79]), .outData_80(wire_con_in_stage3[80]), .outData_81(wire_con_in_stage3[81]), .outData_82(wire_con_in_stage3[82]), .outData_83(wire_con_in_stage3[83]), .outData_84(wire_con_in_stage3[84]), .outData_85(wire_con_in_stage3[85]), .outData_86(wire_con_in_stage3[86]), .outData_87(wire_con_in_stage3[87]), .outData_88(wire_con_in_stage3[88]), .outData_89(wire_con_in_stage3[89]), .outData_90(wire_con_in_stage3[90]), .outData_91(wire_con_in_stage3[91]), .outData_92(wire_con_in_stage3[92]), .outData_93(wire_con_in_stage3[93]), .outData_94(wire_con_in_stage3[94]), .outData_95(wire_con_in_stage3[95]), .outData_96(wire_con_in_stage3[96]), .outData_97(wire_con_in_stage3[97]), .outData_98(wire_con_in_stage3[98]), .outData_99(wire_con_in_stage3[99]), .outData_100(wire_con_in_stage3[100]), .outData_101(wire_con_in_stage3[101]), .outData_102(wire_con_in_stage3[102]), .outData_103(wire_con_in_stage3[103]), .outData_104(wire_con_in_stage3[104]), .outData_105(wire_con_in_stage3[105]), .outData_106(wire_con_in_stage3[106]), .outData_107(wire_con_in_stage3[107]), .outData_108(wire_con_in_stage3[108]), .outData_109(wire_con_in_stage3[109]), .outData_110(wire_con_in_stage3[110]), .outData_111(wire_con_in_stage3[111]), .outData_112(wire_con_in_stage3[112]), .outData_113(wire_con_in_stage3[113]), .outData_114(wire_con_in_stage3[114]), .outData_115(wire_con_in_stage3[115]), .outData_116(wire_con_in_stage3[116]), .outData_117(wire_con_in_stage3[117]), .outData_118(wire_con_in_stage3[118]), .outData_119(wire_con_in_stage3[119]), .outData_120(wire_con_in_stage3[120]), .outData_121(wire_con_in_stage3[121]), .outData_122(wire_con_in_stage3[122]), .outData_123(wire_con_in_stage3[123]), .outData_124(wire_con_in_stage3[124]), .outData_125(wire_con_in_stage3[125]), .outData_126(wire_con_in_stage3[126]), .outData_127(wire_con_in_stage3[127]), .outData_128(wire_con_in_stage3[128]), .outData_129(wire_con_in_stage3[129]), .outData_130(wire_con_in_stage3[130]), .outData_131(wire_con_in_stage3[131]), .outData_132(wire_con_in_stage3[132]), .outData_133(wire_con_in_stage3[133]), .outData_134(wire_con_in_stage3[134]), .outData_135(wire_con_in_stage3[135]), .outData_136(wire_con_in_stage3[136]), .outData_137(wire_con_in_stage3[137]), .outData_138(wire_con_in_stage3[138]), .outData_139(wire_con_in_stage3[139]), .outData_140(wire_con_in_stage3[140]), .outData_141(wire_con_in_stage3[141]), .outData_142(wire_con_in_stage3[142]), .outData_143(wire_con_in_stage3[143]), .outData_144(wire_con_in_stage3[144]), .outData_145(wire_con_in_stage3[145]), .outData_146(wire_con_in_stage3[146]), .outData_147(wire_con_in_stage3[147]), .outData_148(wire_con_in_stage3[148]), .outData_149(wire_con_in_stage3[149]), .outData_150(wire_con_in_stage3[150]), .outData_151(wire_con_in_stage3[151]), .outData_152(wire_con_in_stage3[152]), .outData_153(wire_con_in_stage3[153]), .outData_154(wire_con_in_stage3[154]), .outData_155(wire_con_in_stage3[155]), .outData_156(wire_con_in_stage3[156]), .outData_157(wire_con_in_stage3[157]), .outData_158(wire_con_in_stage3[158]), .outData_159(wire_con_in_stage3[159]), .outData_160(wire_con_in_stage3[160]), .outData_161(wire_con_in_stage3[161]), .outData_162(wire_con_in_stage3[162]), .outData_163(wire_con_in_stage3[163]), .outData_164(wire_con_in_stage3[164]), .outData_165(wire_con_in_stage3[165]), .outData_166(wire_con_in_stage3[166]), .outData_167(wire_con_in_stage3[167]), .outData_168(wire_con_in_stage3[168]), .outData_169(wire_con_in_stage3[169]), .outData_170(wire_con_in_stage3[170]), .outData_171(wire_con_in_stage3[171]), .outData_172(wire_con_in_stage3[172]), .outData_173(wire_con_in_stage3[173]), .outData_174(wire_con_in_stage3[174]), .outData_175(wire_con_in_stage3[175]), .outData_176(wire_con_in_stage3[176]), .outData_177(wire_con_in_stage3[177]), .outData_178(wire_con_in_stage3[178]), .outData_179(wire_con_in_stage3[179]), .outData_180(wire_con_in_stage3[180]), .outData_181(wire_con_in_stage3[181]), .outData_182(wire_con_in_stage3[182]), .outData_183(wire_con_in_stage3[183]), .outData_184(wire_con_in_stage3[184]), .outData_185(wire_con_in_stage3[185]), .outData_186(wire_con_in_stage3[186]), .outData_187(wire_con_in_stage3[187]), .outData_188(wire_con_in_stage3[188]), .outData_189(wire_con_in_stage3[189]), .outData_190(wire_con_in_stage3[190]), .outData_191(wire_con_in_stage3[191]), .outData_192(wire_con_in_stage3[192]), .outData_193(wire_con_in_stage3[193]), .outData_194(wire_con_in_stage3[194]), .outData_195(wire_con_in_stage3[195]), .outData_196(wire_con_in_stage3[196]), .outData_197(wire_con_in_stage3[197]), .outData_198(wire_con_in_stage3[198]), .outData_199(wire_con_in_stage3[199]), .outData_200(wire_con_in_stage3[200]), .outData_201(wire_con_in_stage3[201]), .outData_202(wire_con_in_stage3[202]), .outData_203(wire_con_in_stage3[203]), .outData_204(wire_con_in_stage3[204]), .outData_205(wire_con_in_stage3[205]), .outData_206(wire_con_in_stage3[206]), .outData_207(wire_con_in_stage3[207]), .outData_208(wire_con_in_stage3[208]), .outData_209(wire_con_in_stage3[209]), .outData_210(wire_con_in_stage3[210]), .outData_211(wire_con_in_stage3[211]), .outData_212(wire_con_in_stage3[212]), .outData_213(wire_con_in_stage3[213]), .outData_214(wire_con_in_stage3[214]), .outData_215(wire_con_in_stage3[215]), .outData_216(wire_con_in_stage3[216]), .outData_217(wire_con_in_stage3[217]), .outData_218(wire_con_in_stage3[218]), .outData_219(wire_con_in_stage3[219]), .outData_220(wire_con_in_stage3[220]), .outData_221(wire_con_in_stage3[221]), .outData_222(wire_con_in_stage3[222]), .outData_223(wire_con_in_stage3[223]), .outData_224(wire_con_in_stage3[224]), .outData_225(wire_con_in_stage3[225]), .outData_226(wire_con_in_stage3[226]), .outData_227(wire_con_in_stage3[227]), .outData_228(wire_con_in_stage3[228]), .outData_229(wire_con_in_stage3[229]), .outData_230(wire_con_in_stage3[230]), .outData_231(wire_con_in_stage3[231]), .outData_232(wire_con_in_stage3[232]), .outData_233(wire_con_in_stage3[233]), .outData_234(wire_con_in_stage3[234]), .outData_235(wire_con_in_stage3[235]), .outData_236(wire_con_in_stage3[236]), .outData_237(wire_con_in_stage3[237]), .outData_238(wire_con_in_stage3[238]), .outData_239(wire_con_in_stage3[239]), .outData_240(wire_con_in_stage3[240]), .outData_241(wire_con_in_stage3[241]), .outData_242(wire_con_in_stage3[242]), .outData_243(wire_con_in_stage3[243]), .outData_244(wire_con_in_stage3[244]), .outData_245(wire_con_in_stage3[245]), .outData_246(wire_con_in_stage3[246]), .outData_247(wire_con_in_stage3[247]), .outData_248(wire_con_in_stage3[248]), .outData_249(wire_con_in_stage3[249]), .outData_250(wire_con_in_stage3[250]), .outData_251(wire_con_in_stage3[251]), .outData_252(wire_con_in_stage3[252]), .outData_253(wire_con_in_stage3[253]), .outData_254(wire_con_in_stage3[254]), .outData_255(wire_con_in_stage3[255]), 
        .in_start(in_start_stage3), .out_start(con_in_start_stage3), .ctrl(wire_ctrl_stage3), .clk(clk), .rst(rst));
  
  wireCon_dp256_st3_L wire_stage_3(
        .inData_0(wire_con_in_stage3[0]), .inData_1(wire_con_in_stage3[1]), .inData_2(wire_con_in_stage3[2]), .inData_3(wire_con_in_stage3[3]), .inData_4(wire_con_in_stage3[4]), .inData_5(wire_con_in_stage3[5]), .inData_6(wire_con_in_stage3[6]), .inData_7(wire_con_in_stage3[7]), .inData_8(wire_con_in_stage3[8]), .inData_9(wire_con_in_stage3[9]), .inData_10(wire_con_in_stage3[10]), .inData_11(wire_con_in_stage3[11]), .inData_12(wire_con_in_stage3[12]), .inData_13(wire_con_in_stage3[13]), .inData_14(wire_con_in_stage3[14]), .inData_15(wire_con_in_stage3[15]), .inData_16(wire_con_in_stage3[16]), .inData_17(wire_con_in_stage3[17]), .inData_18(wire_con_in_stage3[18]), .inData_19(wire_con_in_stage3[19]), .inData_20(wire_con_in_stage3[20]), .inData_21(wire_con_in_stage3[21]), .inData_22(wire_con_in_stage3[22]), .inData_23(wire_con_in_stage3[23]), .inData_24(wire_con_in_stage3[24]), .inData_25(wire_con_in_stage3[25]), .inData_26(wire_con_in_stage3[26]), .inData_27(wire_con_in_stage3[27]), .inData_28(wire_con_in_stage3[28]), .inData_29(wire_con_in_stage3[29]), .inData_30(wire_con_in_stage3[30]), .inData_31(wire_con_in_stage3[31]), .inData_32(wire_con_in_stage3[32]), .inData_33(wire_con_in_stage3[33]), .inData_34(wire_con_in_stage3[34]), .inData_35(wire_con_in_stage3[35]), .inData_36(wire_con_in_stage3[36]), .inData_37(wire_con_in_stage3[37]), .inData_38(wire_con_in_stage3[38]), .inData_39(wire_con_in_stage3[39]), .inData_40(wire_con_in_stage3[40]), .inData_41(wire_con_in_stage3[41]), .inData_42(wire_con_in_stage3[42]), .inData_43(wire_con_in_stage3[43]), .inData_44(wire_con_in_stage3[44]), .inData_45(wire_con_in_stage3[45]), .inData_46(wire_con_in_stage3[46]), .inData_47(wire_con_in_stage3[47]), .inData_48(wire_con_in_stage3[48]), .inData_49(wire_con_in_stage3[49]), .inData_50(wire_con_in_stage3[50]), .inData_51(wire_con_in_stage3[51]), .inData_52(wire_con_in_stage3[52]), .inData_53(wire_con_in_stage3[53]), .inData_54(wire_con_in_stage3[54]), .inData_55(wire_con_in_stage3[55]), .inData_56(wire_con_in_stage3[56]), .inData_57(wire_con_in_stage3[57]), .inData_58(wire_con_in_stage3[58]), .inData_59(wire_con_in_stage3[59]), .inData_60(wire_con_in_stage3[60]), .inData_61(wire_con_in_stage3[61]), .inData_62(wire_con_in_stage3[62]), .inData_63(wire_con_in_stage3[63]), .inData_64(wire_con_in_stage3[64]), .inData_65(wire_con_in_stage3[65]), .inData_66(wire_con_in_stage3[66]), .inData_67(wire_con_in_stage3[67]), .inData_68(wire_con_in_stage3[68]), .inData_69(wire_con_in_stage3[69]), .inData_70(wire_con_in_stage3[70]), .inData_71(wire_con_in_stage3[71]), .inData_72(wire_con_in_stage3[72]), .inData_73(wire_con_in_stage3[73]), .inData_74(wire_con_in_stage3[74]), .inData_75(wire_con_in_stage3[75]), .inData_76(wire_con_in_stage3[76]), .inData_77(wire_con_in_stage3[77]), .inData_78(wire_con_in_stage3[78]), .inData_79(wire_con_in_stage3[79]), .inData_80(wire_con_in_stage3[80]), .inData_81(wire_con_in_stage3[81]), .inData_82(wire_con_in_stage3[82]), .inData_83(wire_con_in_stage3[83]), .inData_84(wire_con_in_stage3[84]), .inData_85(wire_con_in_stage3[85]), .inData_86(wire_con_in_stage3[86]), .inData_87(wire_con_in_stage3[87]), .inData_88(wire_con_in_stage3[88]), .inData_89(wire_con_in_stage3[89]), .inData_90(wire_con_in_stage3[90]), .inData_91(wire_con_in_stage3[91]), .inData_92(wire_con_in_stage3[92]), .inData_93(wire_con_in_stage3[93]), .inData_94(wire_con_in_stage3[94]), .inData_95(wire_con_in_stage3[95]), .inData_96(wire_con_in_stage3[96]), .inData_97(wire_con_in_stage3[97]), .inData_98(wire_con_in_stage3[98]), .inData_99(wire_con_in_stage3[99]), .inData_100(wire_con_in_stage3[100]), .inData_101(wire_con_in_stage3[101]), .inData_102(wire_con_in_stage3[102]), .inData_103(wire_con_in_stage3[103]), .inData_104(wire_con_in_stage3[104]), .inData_105(wire_con_in_stage3[105]), .inData_106(wire_con_in_stage3[106]), .inData_107(wire_con_in_stage3[107]), .inData_108(wire_con_in_stage3[108]), .inData_109(wire_con_in_stage3[109]), .inData_110(wire_con_in_stage3[110]), .inData_111(wire_con_in_stage3[111]), .inData_112(wire_con_in_stage3[112]), .inData_113(wire_con_in_stage3[113]), .inData_114(wire_con_in_stage3[114]), .inData_115(wire_con_in_stage3[115]), .inData_116(wire_con_in_stage3[116]), .inData_117(wire_con_in_stage3[117]), .inData_118(wire_con_in_stage3[118]), .inData_119(wire_con_in_stage3[119]), .inData_120(wire_con_in_stage3[120]), .inData_121(wire_con_in_stage3[121]), .inData_122(wire_con_in_stage3[122]), .inData_123(wire_con_in_stage3[123]), .inData_124(wire_con_in_stage3[124]), .inData_125(wire_con_in_stage3[125]), .inData_126(wire_con_in_stage3[126]), .inData_127(wire_con_in_stage3[127]), .inData_128(wire_con_in_stage3[128]), .inData_129(wire_con_in_stage3[129]), .inData_130(wire_con_in_stage3[130]), .inData_131(wire_con_in_stage3[131]), .inData_132(wire_con_in_stage3[132]), .inData_133(wire_con_in_stage3[133]), .inData_134(wire_con_in_stage3[134]), .inData_135(wire_con_in_stage3[135]), .inData_136(wire_con_in_stage3[136]), .inData_137(wire_con_in_stage3[137]), .inData_138(wire_con_in_stage3[138]), .inData_139(wire_con_in_stage3[139]), .inData_140(wire_con_in_stage3[140]), .inData_141(wire_con_in_stage3[141]), .inData_142(wire_con_in_stage3[142]), .inData_143(wire_con_in_stage3[143]), .inData_144(wire_con_in_stage3[144]), .inData_145(wire_con_in_stage3[145]), .inData_146(wire_con_in_stage3[146]), .inData_147(wire_con_in_stage3[147]), .inData_148(wire_con_in_stage3[148]), .inData_149(wire_con_in_stage3[149]), .inData_150(wire_con_in_stage3[150]), .inData_151(wire_con_in_stage3[151]), .inData_152(wire_con_in_stage3[152]), .inData_153(wire_con_in_stage3[153]), .inData_154(wire_con_in_stage3[154]), .inData_155(wire_con_in_stage3[155]), .inData_156(wire_con_in_stage3[156]), .inData_157(wire_con_in_stage3[157]), .inData_158(wire_con_in_stage3[158]), .inData_159(wire_con_in_stage3[159]), .inData_160(wire_con_in_stage3[160]), .inData_161(wire_con_in_stage3[161]), .inData_162(wire_con_in_stage3[162]), .inData_163(wire_con_in_stage3[163]), .inData_164(wire_con_in_stage3[164]), .inData_165(wire_con_in_stage3[165]), .inData_166(wire_con_in_stage3[166]), .inData_167(wire_con_in_stage3[167]), .inData_168(wire_con_in_stage3[168]), .inData_169(wire_con_in_stage3[169]), .inData_170(wire_con_in_stage3[170]), .inData_171(wire_con_in_stage3[171]), .inData_172(wire_con_in_stage3[172]), .inData_173(wire_con_in_stage3[173]), .inData_174(wire_con_in_stage3[174]), .inData_175(wire_con_in_stage3[175]), .inData_176(wire_con_in_stage3[176]), .inData_177(wire_con_in_stage3[177]), .inData_178(wire_con_in_stage3[178]), .inData_179(wire_con_in_stage3[179]), .inData_180(wire_con_in_stage3[180]), .inData_181(wire_con_in_stage3[181]), .inData_182(wire_con_in_stage3[182]), .inData_183(wire_con_in_stage3[183]), .inData_184(wire_con_in_stage3[184]), .inData_185(wire_con_in_stage3[185]), .inData_186(wire_con_in_stage3[186]), .inData_187(wire_con_in_stage3[187]), .inData_188(wire_con_in_stage3[188]), .inData_189(wire_con_in_stage3[189]), .inData_190(wire_con_in_stage3[190]), .inData_191(wire_con_in_stage3[191]), .inData_192(wire_con_in_stage3[192]), .inData_193(wire_con_in_stage3[193]), .inData_194(wire_con_in_stage3[194]), .inData_195(wire_con_in_stage3[195]), .inData_196(wire_con_in_stage3[196]), .inData_197(wire_con_in_stage3[197]), .inData_198(wire_con_in_stage3[198]), .inData_199(wire_con_in_stage3[199]), .inData_200(wire_con_in_stage3[200]), .inData_201(wire_con_in_stage3[201]), .inData_202(wire_con_in_stage3[202]), .inData_203(wire_con_in_stage3[203]), .inData_204(wire_con_in_stage3[204]), .inData_205(wire_con_in_stage3[205]), .inData_206(wire_con_in_stage3[206]), .inData_207(wire_con_in_stage3[207]), .inData_208(wire_con_in_stage3[208]), .inData_209(wire_con_in_stage3[209]), .inData_210(wire_con_in_stage3[210]), .inData_211(wire_con_in_stage3[211]), .inData_212(wire_con_in_stage3[212]), .inData_213(wire_con_in_stage3[213]), .inData_214(wire_con_in_stage3[214]), .inData_215(wire_con_in_stage3[215]), .inData_216(wire_con_in_stage3[216]), .inData_217(wire_con_in_stage3[217]), .inData_218(wire_con_in_stage3[218]), .inData_219(wire_con_in_stage3[219]), .inData_220(wire_con_in_stage3[220]), .inData_221(wire_con_in_stage3[221]), .inData_222(wire_con_in_stage3[222]), .inData_223(wire_con_in_stage3[223]), .inData_224(wire_con_in_stage3[224]), .inData_225(wire_con_in_stage3[225]), .inData_226(wire_con_in_stage3[226]), .inData_227(wire_con_in_stage3[227]), .inData_228(wire_con_in_stage3[228]), .inData_229(wire_con_in_stage3[229]), .inData_230(wire_con_in_stage3[230]), .inData_231(wire_con_in_stage3[231]), .inData_232(wire_con_in_stage3[232]), .inData_233(wire_con_in_stage3[233]), .inData_234(wire_con_in_stage3[234]), .inData_235(wire_con_in_stage3[235]), .inData_236(wire_con_in_stage3[236]), .inData_237(wire_con_in_stage3[237]), .inData_238(wire_con_in_stage3[238]), .inData_239(wire_con_in_stage3[239]), .inData_240(wire_con_in_stage3[240]), .inData_241(wire_con_in_stage3[241]), .inData_242(wire_con_in_stage3[242]), .inData_243(wire_con_in_stage3[243]), .inData_244(wire_con_in_stage3[244]), .inData_245(wire_con_in_stage3[245]), .inData_246(wire_con_in_stage3[246]), .inData_247(wire_con_in_stage3[247]), .inData_248(wire_con_in_stage3[248]), .inData_249(wire_con_in_stage3[249]), .inData_250(wire_con_in_stage3[250]), .inData_251(wire_con_in_stage3[251]), .inData_252(wire_con_in_stage3[252]), .inData_253(wire_con_in_stage3[253]), .inData_254(wire_con_in_stage3[254]), .inData_255(wire_con_in_stage3[255]), 
        .outData_0(wire_con_out_stage3[0]), .outData_1(wire_con_out_stage3[1]), .outData_2(wire_con_out_stage3[2]), .outData_3(wire_con_out_stage3[3]), .outData_4(wire_con_out_stage3[4]), .outData_5(wire_con_out_stage3[5]), .outData_6(wire_con_out_stage3[6]), .outData_7(wire_con_out_stage3[7]), .outData_8(wire_con_out_stage3[8]), .outData_9(wire_con_out_stage3[9]), .outData_10(wire_con_out_stage3[10]), .outData_11(wire_con_out_stage3[11]), .outData_12(wire_con_out_stage3[12]), .outData_13(wire_con_out_stage3[13]), .outData_14(wire_con_out_stage3[14]), .outData_15(wire_con_out_stage3[15]), .outData_16(wire_con_out_stage3[16]), .outData_17(wire_con_out_stage3[17]), .outData_18(wire_con_out_stage3[18]), .outData_19(wire_con_out_stage3[19]), .outData_20(wire_con_out_stage3[20]), .outData_21(wire_con_out_stage3[21]), .outData_22(wire_con_out_stage3[22]), .outData_23(wire_con_out_stage3[23]), .outData_24(wire_con_out_stage3[24]), .outData_25(wire_con_out_stage3[25]), .outData_26(wire_con_out_stage3[26]), .outData_27(wire_con_out_stage3[27]), .outData_28(wire_con_out_stage3[28]), .outData_29(wire_con_out_stage3[29]), .outData_30(wire_con_out_stage3[30]), .outData_31(wire_con_out_stage3[31]), .outData_32(wire_con_out_stage3[32]), .outData_33(wire_con_out_stage3[33]), .outData_34(wire_con_out_stage3[34]), .outData_35(wire_con_out_stage3[35]), .outData_36(wire_con_out_stage3[36]), .outData_37(wire_con_out_stage3[37]), .outData_38(wire_con_out_stage3[38]), .outData_39(wire_con_out_stage3[39]), .outData_40(wire_con_out_stage3[40]), .outData_41(wire_con_out_stage3[41]), .outData_42(wire_con_out_stage3[42]), .outData_43(wire_con_out_stage3[43]), .outData_44(wire_con_out_stage3[44]), .outData_45(wire_con_out_stage3[45]), .outData_46(wire_con_out_stage3[46]), .outData_47(wire_con_out_stage3[47]), .outData_48(wire_con_out_stage3[48]), .outData_49(wire_con_out_stage3[49]), .outData_50(wire_con_out_stage3[50]), .outData_51(wire_con_out_stage3[51]), .outData_52(wire_con_out_stage3[52]), .outData_53(wire_con_out_stage3[53]), .outData_54(wire_con_out_stage3[54]), .outData_55(wire_con_out_stage3[55]), .outData_56(wire_con_out_stage3[56]), .outData_57(wire_con_out_stage3[57]), .outData_58(wire_con_out_stage3[58]), .outData_59(wire_con_out_stage3[59]), .outData_60(wire_con_out_stage3[60]), .outData_61(wire_con_out_stage3[61]), .outData_62(wire_con_out_stage3[62]), .outData_63(wire_con_out_stage3[63]), .outData_64(wire_con_out_stage3[64]), .outData_65(wire_con_out_stage3[65]), .outData_66(wire_con_out_stage3[66]), .outData_67(wire_con_out_stage3[67]), .outData_68(wire_con_out_stage3[68]), .outData_69(wire_con_out_stage3[69]), .outData_70(wire_con_out_stage3[70]), .outData_71(wire_con_out_stage3[71]), .outData_72(wire_con_out_stage3[72]), .outData_73(wire_con_out_stage3[73]), .outData_74(wire_con_out_stage3[74]), .outData_75(wire_con_out_stage3[75]), .outData_76(wire_con_out_stage3[76]), .outData_77(wire_con_out_stage3[77]), .outData_78(wire_con_out_stage3[78]), .outData_79(wire_con_out_stage3[79]), .outData_80(wire_con_out_stage3[80]), .outData_81(wire_con_out_stage3[81]), .outData_82(wire_con_out_stage3[82]), .outData_83(wire_con_out_stage3[83]), .outData_84(wire_con_out_stage3[84]), .outData_85(wire_con_out_stage3[85]), .outData_86(wire_con_out_stage3[86]), .outData_87(wire_con_out_stage3[87]), .outData_88(wire_con_out_stage3[88]), .outData_89(wire_con_out_stage3[89]), .outData_90(wire_con_out_stage3[90]), .outData_91(wire_con_out_stage3[91]), .outData_92(wire_con_out_stage3[92]), .outData_93(wire_con_out_stage3[93]), .outData_94(wire_con_out_stage3[94]), .outData_95(wire_con_out_stage3[95]), .outData_96(wire_con_out_stage3[96]), .outData_97(wire_con_out_stage3[97]), .outData_98(wire_con_out_stage3[98]), .outData_99(wire_con_out_stage3[99]), .outData_100(wire_con_out_stage3[100]), .outData_101(wire_con_out_stage3[101]), .outData_102(wire_con_out_stage3[102]), .outData_103(wire_con_out_stage3[103]), .outData_104(wire_con_out_stage3[104]), .outData_105(wire_con_out_stage3[105]), .outData_106(wire_con_out_stage3[106]), .outData_107(wire_con_out_stage3[107]), .outData_108(wire_con_out_stage3[108]), .outData_109(wire_con_out_stage3[109]), .outData_110(wire_con_out_stage3[110]), .outData_111(wire_con_out_stage3[111]), .outData_112(wire_con_out_stage3[112]), .outData_113(wire_con_out_stage3[113]), .outData_114(wire_con_out_stage3[114]), .outData_115(wire_con_out_stage3[115]), .outData_116(wire_con_out_stage3[116]), .outData_117(wire_con_out_stage3[117]), .outData_118(wire_con_out_stage3[118]), .outData_119(wire_con_out_stage3[119]), .outData_120(wire_con_out_stage3[120]), .outData_121(wire_con_out_stage3[121]), .outData_122(wire_con_out_stage3[122]), .outData_123(wire_con_out_stage3[123]), .outData_124(wire_con_out_stage3[124]), .outData_125(wire_con_out_stage3[125]), .outData_126(wire_con_out_stage3[126]), .outData_127(wire_con_out_stage3[127]), .outData_128(wire_con_out_stage3[128]), .outData_129(wire_con_out_stage3[129]), .outData_130(wire_con_out_stage3[130]), .outData_131(wire_con_out_stage3[131]), .outData_132(wire_con_out_stage3[132]), .outData_133(wire_con_out_stage3[133]), .outData_134(wire_con_out_stage3[134]), .outData_135(wire_con_out_stage3[135]), .outData_136(wire_con_out_stage3[136]), .outData_137(wire_con_out_stage3[137]), .outData_138(wire_con_out_stage3[138]), .outData_139(wire_con_out_stage3[139]), .outData_140(wire_con_out_stage3[140]), .outData_141(wire_con_out_stage3[141]), .outData_142(wire_con_out_stage3[142]), .outData_143(wire_con_out_stage3[143]), .outData_144(wire_con_out_stage3[144]), .outData_145(wire_con_out_stage3[145]), .outData_146(wire_con_out_stage3[146]), .outData_147(wire_con_out_stage3[147]), .outData_148(wire_con_out_stage3[148]), .outData_149(wire_con_out_stage3[149]), .outData_150(wire_con_out_stage3[150]), .outData_151(wire_con_out_stage3[151]), .outData_152(wire_con_out_stage3[152]), .outData_153(wire_con_out_stage3[153]), .outData_154(wire_con_out_stage3[154]), .outData_155(wire_con_out_stage3[155]), .outData_156(wire_con_out_stage3[156]), .outData_157(wire_con_out_stage3[157]), .outData_158(wire_con_out_stage3[158]), .outData_159(wire_con_out_stage3[159]), .outData_160(wire_con_out_stage3[160]), .outData_161(wire_con_out_stage3[161]), .outData_162(wire_con_out_stage3[162]), .outData_163(wire_con_out_stage3[163]), .outData_164(wire_con_out_stage3[164]), .outData_165(wire_con_out_stage3[165]), .outData_166(wire_con_out_stage3[166]), .outData_167(wire_con_out_stage3[167]), .outData_168(wire_con_out_stage3[168]), .outData_169(wire_con_out_stage3[169]), .outData_170(wire_con_out_stage3[170]), .outData_171(wire_con_out_stage3[171]), .outData_172(wire_con_out_stage3[172]), .outData_173(wire_con_out_stage3[173]), .outData_174(wire_con_out_stage3[174]), .outData_175(wire_con_out_stage3[175]), .outData_176(wire_con_out_stage3[176]), .outData_177(wire_con_out_stage3[177]), .outData_178(wire_con_out_stage3[178]), .outData_179(wire_con_out_stage3[179]), .outData_180(wire_con_out_stage3[180]), .outData_181(wire_con_out_stage3[181]), .outData_182(wire_con_out_stage3[182]), .outData_183(wire_con_out_stage3[183]), .outData_184(wire_con_out_stage3[184]), .outData_185(wire_con_out_stage3[185]), .outData_186(wire_con_out_stage3[186]), .outData_187(wire_con_out_stage3[187]), .outData_188(wire_con_out_stage3[188]), .outData_189(wire_con_out_stage3[189]), .outData_190(wire_con_out_stage3[190]), .outData_191(wire_con_out_stage3[191]), .outData_192(wire_con_out_stage3[192]), .outData_193(wire_con_out_stage3[193]), .outData_194(wire_con_out_stage3[194]), .outData_195(wire_con_out_stage3[195]), .outData_196(wire_con_out_stage3[196]), .outData_197(wire_con_out_stage3[197]), .outData_198(wire_con_out_stage3[198]), .outData_199(wire_con_out_stage3[199]), .outData_200(wire_con_out_stage3[200]), .outData_201(wire_con_out_stage3[201]), .outData_202(wire_con_out_stage3[202]), .outData_203(wire_con_out_stage3[203]), .outData_204(wire_con_out_stage3[204]), .outData_205(wire_con_out_stage3[205]), .outData_206(wire_con_out_stage3[206]), .outData_207(wire_con_out_stage3[207]), .outData_208(wire_con_out_stage3[208]), .outData_209(wire_con_out_stage3[209]), .outData_210(wire_con_out_stage3[210]), .outData_211(wire_con_out_stage3[211]), .outData_212(wire_con_out_stage3[212]), .outData_213(wire_con_out_stage3[213]), .outData_214(wire_con_out_stage3[214]), .outData_215(wire_con_out_stage3[215]), .outData_216(wire_con_out_stage3[216]), .outData_217(wire_con_out_stage3[217]), .outData_218(wire_con_out_stage3[218]), .outData_219(wire_con_out_stage3[219]), .outData_220(wire_con_out_stage3[220]), .outData_221(wire_con_out_stage3[221]), .outData_222(wire_con_out_stage3[222]), .outData_223(wire_con_out_stage3[223]), .outData_224(wire_con_out_stage3[224]), .outData_225(wire_con_out_stage3[225]), .outData_226(wire_con_out_stage3[226]), .outData_227(wire_con_out_stage3[227]), .outData_228(wire_con_out_stage3[228]), .outData_229(wire_con_out_stage3[229]), .outData_230(wire_con_out_stage3[230]), .outData_231(wire_con_out_stage3[231]), .outData_232(wire_con_out_stage3[232]), .outData_233(wire_con_out_stage3[233]), .outData_234(wire_con_out_stage3[234]), .outData_235(wire_con_out_stage3[235]), .outData_236(wire_con_out_stage3[236]), .outData_237(wire_con_out_stage3[237]), .outData_238(wire_con_out_stage3[238]), .outData_239(wire_con_out_stage3[239]), .outData_240(wire_con_out_stage3[240]), .outData_241(wire_con_out_stage3[241]), .outData_242(wire_con_out_stage3[242]), .outData_243(wire_con_out_stage3[243]), .outData_244(wire_con_out_stage3[244]), .outData_245(wire_con_out_stage3[245]), .outData_246(wire_con_out_stage3[246]), .outData_247(wire_con_out_stage3[247]), .outData_248(wire_con_out_stage3[248]), .outData_249(wire_con_out_stage3[249]), .outData_250(wire_con_out_stage3[250]), .outData_251(wire_con_out_stage3[251]), .outData_252(wire_con_out_stage3[252]), .outData_253(wire_con_out_stage3[253]), .outData_254(wire_con_out_stage3[254]), .outData_255(wire_con_out_stage3[255]), 
        .in_start(con_in_start_stage3), .out_start(in_start_stage4), .clk(clk), .rst(rst)); 

  
  assign wire_ctrl_stage3[0] = counter_w[4]; 
  assign wire_ctrl_stage3[1] = counter_w[4]; 
  assign wire_ctrl_stage3[2] = counter_w[4]; 
  assign wire_ctrl_stage3[3] = counter_w[4]; 
  assign wire_ctrl_stage3[4] = counter_w[4]; 
  assign wire_ctrl_stage3[5] = counter_w[4]; 
  assign wire_ctrl_stage3[6] = counter_w[4]; 
  assign wire_ctrl_stage3[7] = counter_w[4]; 
  assign wire_ctrl_stage3[8] = counter_w[4]; 
  assign wire_ctrl_stage3[9] = counter_w[4]; 
  assign wire_ctrl_stage3[10] = counter_w[4]; 
  assign wire_ctrl_stage3[11] = counter_w[4]; 
  assign wire_ctrl_stage3[12] = counter_w[4]; 
  assign wire_ctrl_stage3[13] = counter_w[4]; 
  assign wire_ctrl_stage3[14] = counter_w[4]; 
  assign wire_ctrl_stage3[15] = counter_w[4]; 
  assign wire_ctrl_stage3[16] = counter_w[4]; 
  assign wire_ctrl_stage3[17] = counter_w[4]; 
  assign wire_ctrl_stage3[18] = counter_w[4]; 
  assign wire_ctrl_stage3[19] = counter_w[4]; 
  assign wire_ctrl_stage3[20] = counter_w[4]; 
  assign wire_ctrl_stage3[21] = counter_w[4]; 
  assign wire_ctrl_stage3[22] = counter_w[4]; 
  assign wire_ctrl_stage3[23] = counter_w[4]; 
  assign wire_ctrl_stage3[24] = counter_w[4]; 
  assign wire_ctrl_stage3[25] = counter_w[4]; 
  assign wire_ctrl_stage3[26] = counter_w[4]; 
  assign wire_ctrl_stage3[27] = counter_w[4]; 
  assign wire_ctrl_stage3[28] = counter_w[4]; 
  assign wire_ctrl_stage3[29] = counter_w[4]; 
  assign wire_ctrl_stage3[30] = counter_w[4]; 
  assign wire_ctrl_stage3[31] = counter_w[4]; 
  assign wire_ctrl_stage3[32] = counter_w[4]; 
  assign wire_ctrl_stage3[33] = counter_w[4]; 
  assign wire_ctrl_stage3[34] = counter_w[4]; 
  assign wire_ctrl_stage3[35] = counter_w[4]; 
  assign wire_ctrl_stage3[36] = counter_w[4]; 
  assign wire_ctrl_stage3[37] = counter_w[4]; 
  assign wire_ctrl_stage3[38] = counter_w[4]; 
  assign wire_ctrl_stage3[39] = counter_w[4]; 
  assign wire_ctrl_stage3[40] = counter_w[4]; 
  assign wire_ctrl_stage3[41] = counter_w[4]; 
  assign wire_ctrl_stage3[42] = counter_w[4]; 
  assign wire_ctrl_stage3[43] = counter_w[4]; 
  assign wire_ctrl_stage3[44] = counter_w[4]; 
  assign wire_ctrl_stage3[45] = counter_w[4]; 
  assign wire_ctrl_stage3[46] = counter_w[4]; 
  assign wire_ctrl_stage3[47] = counter_w[4]; 
  assign wire_ctrl_stage3[48] = counter_w[4]; 
  assign wire_ctrl_stage3[49] = counter_w[4]; 
  assign wire_ctrl_stage3[50] = counter_w[4]; 
  assign wire_ctrl_stage3[51] = counter_w[4]; 
  assign wire_ctrl_stage3[52] = counter_w[4]; 
  assign wire_ctrl_stage3[53] = counter_w[4]; 
  assign wire_ctrl_stage3[54] = counter_w[4]; 
  assign wire_ctrl_stage3[55] = counter_w[4]; 
  assign wire_ctrl_stage3[56] = counter_w[4]; 
  assign wire_ctrl_stage3[57] = counter_w[4]; 
  assign wire_ctrl_stage3[58] = counter_w[4]; 
  assign wire_ctrl_stage3[59] = counter_w[4]; 
  assign wire_ctrl_stage3[60] = counter_w[4]; 
  assign wire_ctrl_stage3[61] = counter_w[4]; 
  assign wire_ctrl_stage3[62] = counter_w[4]; 
  assign wire_ctrl_stage3[63] = counter_w[4]; 
  assign wire_ctrl_stage3[64] = counter_w[4]; 
  assign wire_ctrl_stage3[65] = counter_w[4]; 
  assign wire_ctrl_stage3[66] = counter_w[4]; 
  assign wire_ctrl_stage3[67] = counter_w[4]; 
  assign wire_ctrl_stage3[68] = counter_w[4]; 
  assign wire_ctrl_stage3[69] = counter_w[4]; 
  assign wire_ctrl_stage3[70] = counter_w[4]; 
  assign wire_ctrl_stage3[71] = counter_w[4]; 
  assign wire_ctrl_stage3[72] = counter_w[4]; 
  assign wire_ctrl_stage3[73] = counter_w[4]; 
  assign wire_ctrl_stage3[74] = counter_w[4]; 
  assign wire_ctrl_stage3[75] = counter_w[4]; 
  assign wire_ctrl_stage3[76] = counter_w[4]; 
  assign wire_ctrl_stage3[77] = counter_w[4]; 
  assign wire_ctrl_stage3[78] = counter_w[4]; 
  assign wire_ctrl_stage3[79] = counter_w[4]; 
  assign wire_ctrl_stage3[80] = counter_w[4]; 
  assign wire_ctrl_stage3[81] = counter_w[4]; 
  assign wire_ctrl_stage3[82] = counter_w[4]; 
  assign wire_ctrl_stage3[83] = counter_w[4]; 
  assign wire_ctrl_stage3[84] = counter_w[4]; 
  assign wire_ctrl_stage3[85] = counter_w[4]; 
  assign wire_ctrl_stage3[86] = counter_w[4]; 
  assign wire_ctrl_stage3[87] = counter_w[4]; 
  assign wire_ctrl_stage3[88] = counter_w[4]; 
  assign wire_ctrl_stage3[89] = counter_w[4]; 
  assign wire_ctrl_stage3[90] = counter_w[4]; 
  assign wire_ctrl_stage3[91] = counter_w[4]; 
  assign wire_ctrl_stage3[92] = counter_w[4]; 
  assign wire_ctrl_stage3[93] = counter_w[4]; 
  assign wire_ctrl_stage3[94] = counter_w[4]; 
  assign wire_ctrl_stage3[95] = counter_w[4]; 
  assign wire_ctrl_stage3[96] = counter_w[4]; 
  assign wire_ctrl_stage3[97] = counter_w[4]; 
  assign wire_ctrl_stage3[98] = counter_w[4]; 
  assign wire_ctrl_stage3[99] = counter_w[4]; 
  assign wire_ctrl_stage3[100] = counter_w[4]; 
  assign wire_ctrl_stage3[101] = counter_w[4]; 
  assign wire_ctrl_stage3[102] = counter_w[4]; 
  assign wire_ctrl_stage3[103] = counter_w[4]; 
  assign wire_ctrl_stage3[104] = counter_w[4]; 
  assign wire_ctrl_stage3[105] = counter_w[4]; 
  assign wire_ctrl_stage3[106] = counter_w[4]; 
  assign wire_ctrl_stage3[107] = counter_w[4]; 
  assign wire_ctrl_stage3[108] = counter_w[4]; 
  assign wire_ctrl_stage3[109] = counter_w[4]; 
  assign wire_ctrl_stage3[110] = counter_w[4]; 
  assign wire_ctrl_stage3[111] = counter_w[4]; 
  assign wire_ctrl_stage3[112] = counter_w[4]; 
  assign wire_ctrl_stage3[113] = counter_w[4]; 
  assign wire_ctrl_stage3[114] = counter_w[4]; 
  assign wire_ctrl_stage3[115] = counter_w[4]; 
  assign wire_ctrl_stage3[116] = counter_w[4]; 
  assign wire_ctrl_stage3[117] = counter_w[4]; 
  assign wire_ctrl_stage3[118] = counter_w[4]; 
  assign wire_ctrl_stage3[119] = counter_w[4]; 
  assign wire_ctrl_stage3[120] = counter_w[4]; 
  assign wire_ctrl_stage3[121] = counter_w[4]; 
  assign wire_ctrl_stage3[122] = counter_w[4]; 
  assign wire_ctrl_stage3[123] = counter_w[4]; 
  assign wire_ctrl_stage3[124] = counter_w[4]; 
  assign wire_ctrl_stage3[125] = counter_w[4]; 
  assign wire_ctrl_stage3[126] = counter_w[4]; 
  assign wire_ctrl_stage3[127] = counter_w[4]; 
  wire [DATA_WIDTH-1:0] wire_con_in_stage4[255:0];
  wire [DATA_WIDTH-1:0] wire_con_out_stage4[255:0];
  wire [127:0] wire_ctrl_stage4;

  switches_stage_st4_0_L switch_stage_4(
        .inData_0(wire_con_out_stage3[0]), .inData_1(wire_con_out_stage3[1]), .inData_2(wire_con_out_stage3[2]), .inData_3(wire_con_out_stage3[3]), .inData_4(wire_con_out_stage3[4]), .inData_5(wire_con_out_stage3[5]), .inData_6(wire_con_out_stage3[6]), .inData_7(wire_con_out_stage3[7]), .inData_8(wire_con_out_stage3[8]), .inData_9(wire_con_out_stage3[9]), .inData_10(wire_con_out_stage3[10]), .inData_11(wire_con_out_stage3[11]), .inData_12(wire_con_out_stage3[12]), .inData_13(wire_con_out_stage3[13]), .inData_14(wire_con_out_stage3[14]), .inData_15(wire_con_out_stage3[15]), .inData_16(wire_con_out_stage3[16]), .inData_17(wire_con_out_stage3[17]), .inData_18(wire_con_out_stage3[18]), .inData_19(wire_con_out_stage3[19]), .inData_20(wire_con_out_stage3[20]), .inData_21(wire_con_out_stage3[21]), .inData_22(wire_con_out_stage3[22]), .inData_23(wire_con_out_stage3[23]), .inData_24(wire_con_out_stage3[24]), .inData_25(wire_con_out_stage3[25]), .inData_26(wire_con_out_stage3[26]), .inData_27(wire_con_out_stage3[27]), .inData_28(wire_con_out_stage3[28]), .inData_29(wire_con_out_stage3[29]), .inData_30(wire_con_out_stage3[30]), .inData_31(wire_con_out_stage3[31]), .inData_32(wire_con_out_stage3[32]), .inData_33(wire_con_out_stage3[33]), .inData_34(wire_con_out_stage3[34]), .inData_35(wire_con_out_stage3[35]), .inData_36(wire_con_out_stage3[36]), .inData_37(wire_con_out_stage3[37]), .inData_38(wire_con_out_stage3[38]), .inData_39(wire_con_out_stage3[39]), .inData_40(wire_con_out_stage3[40]), .inData_41(wire_con_out_stage3[41]), .inData_42(wire_con_out_stage3[42]), .inData_43(wire_con_out_stage3[43]), .inData_44(wire_con_out_stage3[44]), .inData_45(wire_con_out_stage3[45]), .inData_46(wire_con_out_stage3[46]), .inData_47(wire_con_out_stage3[47]), .inData_48(wire_con_out_stage3[48]), .inData_49(wire_con_out_stage3[49]), .inData_50(wire_con_out_stage3[50]), .inData_51(wire_con_out_stage3[51]), .inData_52(wire_con_out_stage3[52]), .inData_53(wire_con_out_stage3[53]), .inData_54(wire_con_out_stage3[54]), .inData_55(wire_con_out_stage3[55]), .inData_56(wire_con_out_stage3[56]), .inData_57(wire_con_out_stage3[57]), .inData_58(wire_con_out_stage3[58]), .inData_59(wire_con_out_stage3[59]), .inData_60(wire_con_out_stage3[60]), .inData_61(wire_con_out_stage3[61]), .inData_62(wire_con_out_stage3[62]), .inData_63(wire_con_out_stage3[63]), .inData_64(wire_con_out_stage3[64]), .inData_65(wire_con_out_stage3[65]), .inData_66(wire_con_out_stage3[66]), .inData_67(wire_con_out_stage3[67]), .inData_68(wire_con_out_stage3[68]), .inData_69(wire_con_out_stage3[69]), .inData_70(wire_con_out_stage3[70]), .inData_71(wire_con_out_stage3[71]), .inData_72(wire_con_out_stage3[72]), .inData_73(wire_con_out_stage3[73]), .inData_74(wire_con_out_stage3[74]), .inData_75(wire_con_out_stage3[75]), .inData_76(wire_con_out_stage3[76]), .inData_77(wire_con_out_stage3[77]), .inData_78(wire_con_out_stage3[78]), .inData_79(wire_con_out_stage3[79]), .inData_80(wire_con_out_stage3[80]), .inData_81(wire_con_out_stage3[81]), .inData_82(wire_con_out_stage3[82]), .inData_83(wire_con_out_stage3[83]), .inData_84(wire_con_out_stage3[84]), .inData_85(wire_con_out_stage3[85]), .inData_86(wire_con_out_stage3[86]), .inData_87(wire_con_out_stage3[87]), .inData_88(wire_con_out_stage3[88]), .inData_89(wire_con_out_stage3[89]), .inData_90(wire_con_out_stage3[90]), .inData_91(wire_con_out_stage3[91]), .inData_92(wire_con_out_stage3[92]), .inData_93(wire_con_out_stage3[93]), .inData_94(wire_con_out_stage3[94]), .inData_95(wire_con_out_stage3[95]), .inData_96(wire_con_out_stage3[96]), .inData_97(wire_con_out_stage3[97]), .inData_98(wire_con_out_stage3[98]), .inData_99(wire_con_out_stage3[99]), .inData_100(wire_con_out_stage3[100]), .inData_101(wire_con_out_stage3[101]), .inData_102(wire_con_out_stage3[102]), .inData_103(wire_con_out_stage3[103]), .inData_104(wire_con_out_stage3[104]), .inData_105(wire_con_out_stage3[105]), .inData_106(wire_con_out_stage3[106]), .inData_107(wire_con_out_stage3[107]), .inData_108(wire_con_out_stage3[108]), .inData_109(wire_con_out_stage3[109]), .inData_110(wire_con_out_stage3[110]), .inData_111(wire_con_out_stage3[111]), .inData_112(wire_con_out_stage3[112]), .inData_113(wire_con_out_stage3[113]), .inData_114(wire_con_out_stage3[114]), .inData_115(wire_con_out_stage3[115]), .inData_116(wire_con_out_stage3[116]), .inData_117(wire_con_out_stage3[117]), .inData_118(wire_con_out_stage3[118]), .inData_119(wire_con_out_stage3[119]), .inData_120(wire_con_out_stage3[120]), .inData_121(wire_con_out_stage3[121]), .inData_122(wire_con_out_stage3[122]), .inData_123(wire_con_out_stage3[123]), .inData_124(wire_con_out_stage3[124]), .inData_125(wire_con_out_stage3[125]), .inData_126(wire_con_out_stage3[126]), .inData_127(wire_con_out_stage3[127]), .inData_128(wire_con_out_stage3[128]), .inData_129(wire_con_out_stage3[129]), .inData_130(wire_con_out_stage3[130]), .inData_131(wire_con_out_stage3[131]), .inData_132(wire_con_out_stage3[132]), .inData_133(wire_con_out_stage3[133]), .inData_134(wire_con_out_stage3[134]), .inData_135(wire_con_out_stage3[135]), .inData_136(wire_con_out_stage3[136]), .inData_137(wire_con_out_stage3[137]), .inData_138(wire_con_out_stage3[138]), .inData_139(wire_con_out_stage3[139]), .inData_140(wire_con_out_stage3[140]), .inData_141(wire_con_out_stage3[141]), .inData_142(wire_con_out_stage3[142]), .inData_143(wire_con_out_stage3[143]), .inData_144(wire_con_out_stage3[144]), .inData_145(wire_con_out_stage3[145]), .inData_146(wire_con_out_stage3[146]), .inData_147(wire_con_out_stage3[147]), .inData_148(wire_con_out_stage3[148]), .inData_149(wire_con_out_stage3[149]), .inData_150(wire_con_out_stage3[150]), .inData_151(wire_con_out_stage3[151]), .inData_152(wire_con_out_stage3[152]), .inData_153(wire_con_out_stage3[153]), .inData_154(wire_con_out_stage3[154]), .inData_155(wire_con_out_stage3[155]), .inData_156(wire_con_out_stage3[156]), .inData_157(wire_con_out_stage3[157]), .inData_158(wire_con_out_stage3[158]), .inData_159(wire_con_out_stage3[159]), .inData_160(wire_con_out_stage3[160]), .inData_161(wire_con_out_stage3[161]), .inData_162(wire_con_out_stage3[162]), .inData_163(wire_con_out_stage3[163]), .inData_164(wire_con_out_stage3[164]), .inData_165(wire_con_out_stage3[165]), .inData_166(wire_con_out_stage3[166]), .inData_167(wire_con_out_stage3[167]), .inData_168(wire_con_out_stage3[168]), .inData_169(wire_con_out_stage3[169]), .inData_170(wire_con_out_stage3[170]), .inData_171(wire_con_out_stage3[171]), .inData_172(wire_con_out_stage3[172]), .inData_173(wire_con_out_stage3[173]), .inData_174(wire_con_out_stage3[174]), .inData_175(wire_con_out_stage3[175]), .inData_176(wire_con_out_stage3[176]), .inData_177(wire_con_out_stage3[177]), .inData_178(wire_con_out_stage3[178]), .inData_179(wire_con_out_stage3[179]), .inData_180(wire_con_out_stage3[180]), .inData_181(wire_con_out_stage3[181]), .inData_182(wire_con_out_stage3[182]), .inData_183(wire_con_out_stage3[183]), .inData_184(wire_con_out_stage3[184]), .inData_185(wire_con_out_stage3[185]), .inData_186(wire_con_out_stage3[186]), .inData_187(wire_con_out_stage3[187]), .inData_188(wire_con_out_stage3[188]), .inData_189(wire_con_out_stage3[189]), .inData_190(wire_con_out_stage3[190]), .inData_191(wire_con_out_stage3[191]), .inData_192(wire_con_out_stage3[192]), .inData_193(wire_con_out_stage3[193]), .inData_194(wire_con_out_stage3[194]), .inData_195(wire_con_out_stage3[195]), .inData_196(wire_con_out_stage3[196]), .inData_197(wire_con_out_stage3[197]), .inData_198(wire_con_out_stage3[198]), .inData_199(wire_con_out_stage3[199]), .inData_200(wire_con_out_stage3[200]), .inData_201(wire_con_out_stage3[201]), .inData_202(wire_con_out_stage3[202]), .inData_203(wire_con_out_stage3[203]), .inData_204(wire_con_out_stage3[204]), .inData_205(wire_con_out_stage3[205]), .inData_206(wire_con_out_stage3[206]), .inData_207(wire_con_out_stage3[207]), .inData_208(wire_con_out_stage3[208]), .inData_209(wire_con_out_stage3[209]), .inData_210(wire_con_out_stage3[210]), .inData_211(wire_con_out_stage3[211]), .inData_212(wire_con_out_stage3[212]), .inData_213(wire_con_out_stage3[213]), .inData_214(wire_con_out_stage3[214]), .inData_215(wire_con_out_stage3[215]), .inData_216(wire_con_out_stage3[216]), .inData_217(wire_con_out_stage3[217]), .inData_218(wire_con_out_stage3[218]), .inData_219(wire_con_out_stage3[219]), .inData_220(wire_con_out_stage3[220]), .inData_221(wire_con_out_stage3[221]), .inData_222(wire_con_out_stage3[222]), .inData_223(wire_con_out_stage3[223]), .inData_224(wire_con_out_stage3[224]), .inData_225(wire_con_out_stage3[225]), .inData_226(wire_con_out_stage3[226]), .inData_227(wire_con_out_stage3[227]), .inData_228(wire_con_out_stage3[228]), .inData_229(wire_con_out_stage3[229]), .inData_230(wire_con_out_stage3[230]), .inData_231(wire_con_out_stage3[231]), .inData_232(wire_con_out_stage3[232]), .inData_233(wire_con_out_stage3[233]), .inData_234(wire_con_out_stage3[234]), .inData_235(wire_con_out_stage3[235]), .inData_236(wire_con_out_stage3[236]), .inData_237(wire_con_out_stage3[237]), .inData_238(wire_con_out_stage3[238]), .inData_239(wire_con_out_stage3[239]), .inData_240(wire_con_out_stage3[240]), .inData_241(wire_con_out_stage3[241]), .inData_242(wire_con_out_stage3[242]), .inData_243(wire_con_out_stage3[243]), .inData_244(wire_con_out_stage3[244]), .inData_245(wire_con_out_stage3[245]), .inData_246(wire_con_out_stage3[246]), .inData_247(wire_con_out_stage3[247]), .inData_248(wire_con_out_stage3[248]), .inData_249(wire_con_out_stage3[249]), .inData_250(wire_con_out_stage3[250]), .inData_251(wire_con_out_stage3[251]), .inData_252(wire_con_out_stage3[252]), .inData_253(wire_con_out_stage3[253]), .inData_254(wire_con_out_stage3[254]), .inData_255(wire_con_out_stage3[255]), 
        .outData_0(wire_con_in_stage4[0]), .outData_1(wire_con_in_stage4[1]), .outData_2(wire_con_in_stage4[2]), .outData_3(wire_con_in_stage4[3]), .outData_4(wire_con_in_stage4[4]), .outData_5(wire_con_in_stage4[5]), .outData_6(wire_con_in_stage4[6]), .outData_7(wire_con_in_stage4[7]), .outData_8(wire_con_in_stage4[8]), .outData_9(wire_con_in_stage4[9]), .outData_10(wire_con_in_stage4[10]), .outData_11(wire_con_in_stage4[11]), .outData_12(wire_con_in_stage4[12]), .outData_13(wire_con_in_stage4[13]), .outData_14(wire_con_in_stage4[14]), .outData_15(wire_con_in_stage4[15]), .outData_16(wire_con_in_stage4[16]), .outData_17(wire_con_in_stage4[17]), .outData_18(wire_con_in_stage4[18]), .outData_19(wire_con_in_stage4[19]), .outData_20(wire_con_in_stage4[20]), .outData_21(wire_con_in_stage4[21]), .outData_22(wire_con_in_stage4[22]), .outData_23(wire_con_in_stage4[23]), .outData_24(wire_con_in_stage4[24]), .outData_25(wire_con_in_stage4[25]), .outData_26(wire_con_in_stage4[26]), .outData_27(wire_con_in_stage4[27]), .outData_28(wire_con_in_stage4[28]), .outData_29(wire_con_in_stage4[29]), .outData_30(wire_con_in_stage4[30]), .outData_31(wire_con_in_stage4[31]), .outData_32(wire_con_in_stage4[32]), .outData_33(wire_con_in_stage4[33]), .outData_34(wire_con_in_stage4[34]), .outData_35(wire_con_in_stage4[35]), .outData_36(wire_con_in_stage4[36]), .outData_37(wire_con_in_stage4[37]), .outData_38(wire_con_in_stage4[38]), .outData_39(wire_con_in_stage4[39]), .outData_40(wire_con_in_stage4[40]), .outData_41(wire_con_in_stage4[41]), .outData_42(wire_con_in_stage4[42]), .outData_43(wire_con_in_stage4[43]), .outData_44(wire_con_in_stage4[44]), .outData_45(wire_con_in_stage4[45]), .outData_46(wire_con_in_stage4[46]), .outData_47(wire_con_in_stage4[47]), .outData_48(wire_con_in_stage4[48]), .outData_49(wire_con_in_stage4[49]), .outData_50(wire_con_in_stage4[50]), .outData_51(wire_con_in_stage4[51]), .outData_52(wire_con_in_stage4[52]), .outData_53(wire_con_in_stage4[53]), .outData_54(wire_con_in_stage4[54]), .outData_55(wire_con_in_stage4[55]), .outData_56(wire_con_in_stage4[56]), .outData_57(wire_con_in_stage4[57]), .outData_58(wire_con_in_stage4[58]), .outData_59(wire_con_in_stage4[59]), .outData_60(wire_con_in_stage4[60]), .outData_61(wire_con_in_stage4[61]), .outData_62(wire_con_in_stage4[62]), .outData_63(wire_con_in_stage4[63]), .outData_64(wire_con_in_stage4[64]), .outData_65(wire_con_in_stage4[65]), .outData_66(wire_con_in_stage4[66]), .outData_67(wire_con_in_stage4[67]), .outData_68(wire_con_in_stage4[68]), .outData_69(wire_con_in_stage4[69]), .outData_70(wire_con_in_stage4[70]), .outData_71(wire_con_in_stage4[71]), .outData_72(wire_con_in_stage4[72]), .outData_73(wire_con_in_stage4[73]), .outData_74(wire_con_in_stage4[74]), .outData_75(wire_con_in_stage4[75]), .outData_76(wire_con_in_stage4[76]), .outData_77(wire_con_in_stage4[77]), .outData_78(wire_con_in_stage4[78]), .outData_79(wire_con_in_stage4[79]), .outData_80(wire_con_in_stage4[80]), .outData_81(wire_con_in_stage4[81]), .outData_82(wire_con_in_stage4[82]), .outData_83(wire_con_in_stage4[83]), .outData_84(wire_con_in_stage4[84]), .outData_85(wire_con_in_stage4[85]), .outData_86(wire_con_in_stage4[86]), .outData_87(wire_con_in_stage4[87]), .outData_88(wire_con_in_stage4[88]), .outData_89(wire_con_in_stage4[89]), .outData_90(wire_con_in_stage4[90]), .outData_91(wire_con_in_stage4[91]), .outData_92(wire_con_in_stage4[92]), .outData_93(wire_con_in_stage4[93]), .outData_94(wire_con_in_stage4[94]), .outData_95(wire_con_in_stage4[95]), .outData_96(wire_con_in_stage4[96]), .outData_97(wire_con_in_stage4[97]), .outData_98(wire_con_in_stage4[98]), .outData_99(wire_con_in_stage4[99]), .outData_100(wire_con_in_stage4[100]), .outData_101(wire_con_in_stage4[101]), .outData_102(wire_con_in_stage4[102]), .outData_103(wire_con_in_stage4[103]), .outData_104(wire_con_in_stage4[104]), .outData_105(wire_con_in_stage4[105]), .outData_106(wire_con_in_stage4[106]), .outData_107(wire_con_in_stage4[107]), .outData_108(wire_con_in_stage4[108]), .outData_109(wire_con_in_stage4[109]), .outData_110(wire_con_in_stage4[110]), .outData_111(wire_con_in_stage4[111]), .outData_112(wire_con_in_stage4[112]), .outData_113(wire_con_in_stage4[113]), .outData_114(wire_con_in_stage4[114]), .outData_115(wire_con_in_stage4[115]), .outData_116(wire_con_in_stage4[116]), .outData_117(wire_con_in_stage4[117]), .outData_118(wire_con_in_stage4[118]), .outData_119(wire_con_in_stage4[119]), .outData_120(wire_con_in_stage4[120]), .outData_121(wire_con_in_stage4[121]), .outData_122(wire_con_in_stage4[122]), .outData_123(wire_con_in_stage4[123]), .outData_124(wire_con_in_stage4[124]), .outData_125(wire_con_in_stage4[125]), .outData_126(wire_con_in_stage4[126]), .outData_127(wire_con_in_stage4[127]), .outData_128(wire_con_in_stage4[128]), .outData_129(wire_con_in_stage4[129]), .outData_130(wire_con_in_stage4[130]), .outData_131(wire_con_in_stage4[131]), .outData_132(wire_con_in_stage4[132]), .outData_133(wire_con_in_stage4[133]), .outData_134(wire_con_in_stage4[134]), .outData_135(wire_con_in_stage4[135]), .outData_136(wire_con_in_stage4[136]), .outData_137(wire_con_in_stage4[137]), .outData_138(wire_con_in_stage4[138]), .outData_139(wire_con_in_stage4[139]), .outData_140(wire_con_in_stage4[140]), .outData_141(wire_con_in_stage4[141]), .outData_142(wire_con_in_stage4[142]), .outData_143(wire_con_in_stage4[143]), .outData_144(wire_con_in_stage4[144]), .outData_145(wire_con_in_stage4[145]), .outData_146(wire_con_in_stage4[146]), .outData_147(wire_con_in_stage4[147]), .outData_148(wire_con_in_stage4[148]), .outData_149(wire_con_in_stage4[149]), .outData_150(wire_con_in_stage4[150]), .outData_151(wire_con_in_stage4[151]), .outData_152(wire_con_in_stage4[152]), .outData_153(wire_con_in_stage4[153]), .outData_154(wire_con_in_stage4[154]), .outData_155(wire_con_in_stage4[155]), .outData_156(wire_con_in_stage4[156]), .outData_157(wire_con_in_stage4[157]), .outData_158(wire_con_in_stage4[158]), .outData_159(wire_con_in_stage4[159]), .outData_160(wire_con_in_stage4[160]), .outData_161(wire_con_in_stage4[161]), .outData_162(wire_con_in_stage4[162]), .outData_163(wire_con_in_stage4[163]), .outData_164(wire_con_in_stage4[164]), .outData_165(wire_con_in_stage4[165]), .outData_166(wire_con_in_stage4[166]), .outData_167(wire_con_in_stage4[167]), .outData_168(wire_con_in_stage4[168]), .outData_169(wire_con_in_stage4[169]), .outData_170(wire_con_in_stage4[170]), .outData_171(wire_con_in_stage4[171]), .outData_172(wire_con_in_stage4[172]), .outData_173(wire_con_in_stage4[173]), .outData_174(wire_con_in_stage4[174]), .outData_175(wire_con_in_stage4[175]), .outData_176(wire_con_in_stage4[176]), .outData_177(wire_con_in_stage4[177]), .outData_178(wire_con_in_stage4[178]), .outData_179(wire_con_in_stage4[179]), .outData_180(wire_con_in_stage4[180]), .outData_181(wire_con_in_stage4[181]), .outData_182(wire_con_in_stage4[182]), .outData_183(wire_con_in_stage4[183]), .outData_184(wire_con_in_stage4[184]), .outData_185(wire_con_in_stage4[185]), .outData_186(wire_con_in_stage4[186]), .outData_187(wire_con_in_stage4[187]), .outData_188(wire_con_in_stage4[188]), .outData_189(wire_con_in_stage4[189]), .outData_190(wire_con_in_stage4[190]), .outData_191(wire_con_in_stage4[191]), .outData_192(wire_con_in_stage4[192]), .outData_193(wire_con_in_stage4[193]), .outData_194(wire_con_in_stage4[194]), .outData_195(wire_con_in_stage4[195]), .outData_196(wire_con_in_stage4[196]), .outData_197(wire_con_in_stage4[197]), .outData_198(wire_con_in_stage4[198]), .outData_199(wire_con_in_stage4[199]), .outData_200(wire_con_in_stage4[200]), .outData_201(wire_con_in_stage4[201]), .outData_202(wire_con_in_stage4[202]), .outData_203(wire_con_in_stage4[203]), .outData_204(wire_con_in_stage4[204]), .outData_205(wire_con_in_stage4[205]), .outData_206(wire_con_in_stage4[206]), .outData_207(wire_con_in_stage4[207]), .outData_208(wire_con_in_stage4[208]), .outData_209(wire_con_in_stage4[209]), .outData_210(wire_con_in_stage4[210]), .outData_211(wire_con_in_stage4[211]), .outData_212(wire_con_in_stage4[212]), .outData_213(wire_con_in_stage4[213]), .outData_214(wire_con_in_stage4[214]), .outData_215(wire_con_in_stage4[215]), .outData_216(wire_con_in_stage4[216]), .outData_217(wire_con_in_stage4[217]), .outData_218(wire_con_in_stage4[218]), .outData_219(wire_con_in_stage4[219]), .outData_220(wire_con_in_stage4[220]), .outData_221(wire_con_in_stage4[221]), .outData_222(wire_con_in_stage4[222]), .outData_223(wire_con_in_stage4[223]), .outData_224(wire_con_in_stage4[224]), .outData_225(wire_con_in_stage4[225]), .outData_226(wire_con_in_stage4[226]), .outData_227(wire_con_in_stage4[227]), .outData_228(wire_con_in_stage4[228]), .outData_229(wire_con_in_stage4[229]), .outData_230(wire_con_in_stage4[230]), .outData_231(wire_con_in_stage4[231]), .outData_232(wire_con_in_stage4[232]), .outData_233(wire_con_in_stage4[233]), .outData_234(wire_con_in_stage4[234]), .outData_235(wire_con_in_stage4[235]), .outData_236(wire_con_in_stage4[236]), .outData_237(wire_con_in_stage4[237]), .outData_238(wire_con_in_stage4[238]), .outData_239(wire_con_in_stage4[239]), .outData_240(wire_con_in_stage4[240]), .outData_241(wire_con_in_stage4[241]), .outData_242(wire_con_in_stage4[242]), .outData_243(wire_con_in_stage4[243]), .outData_244(wire_con_in_stage4[244]), .outData_245(wire_con_in_stage4[245]), .outData_246(wire_con_in_stage4[246]), .outData_247(wire_con_in_stage4[247]), .outData_248(wire_con_in_stage4[248]), .outData_249(wire_con_in_stage4[249]), .outData_250(wire_con_in_stage4[250]), .outData_251(wire_con_in_stage4[251]), .outData_252(wire_con_in_stage4[252]), .outData_253(wire_con_in_stage4[253]), .outData_254(wire_con_in_stage4[254]), .outData_255(wire_con_in_stage4[255]), 
        .in_start(in_start_stage4), .out_start(con_in_start_stage4), .ctrl(wire_ctrl_stage4), .clk(clk), .rst(rst));
  
  wireCon_dp256_st4_L wire_stage_4(
        .inData_0(wire_con_in_stage4[0]), .inData_1(wire_con_in_stage4[1]), .inData_2(wire_con_in_stage4[2]), .inData_3(wire_con_in_stage4[3]), .inData_4(wire_con_in_stage4[4]), .inData_5(wire_con_in_stage4[5]), .inData_6(wire_con_in_stage4[6]), .inData_7(wire_con_in_stage4[7]), .inData_8(wire_con_in_stage4[8]), .inData_9(wire_con_in_stage4[9]), .inData_10(wire_con_in_stage4[10]), .inData_11(wire_con_in_stage4[11]), .inData_12(wire_con_in_stage4[12]), .inData_13(wire_con_in_stage4[13]), .inData_14(wire_con_in_stage4[14]), .inData_15(wire_con_in_stage4[15]), .inData_16(wire_con_in_stage4[16]), .inData_17(wire_con_in_stage4[17]), .inData_18(wire_con_in_stage4[18]), .inData_19(wire_con_in_stage4[19]), .inData_20(wire_con_in_stage4[20]), .inData_21(wire_con_in_stage4[21]), .inData_22(wire_con_in_stage4[22]), .inData_23(wire_con_in_stage4[23]), .inData_24(wire_con_in_stage4[24]), .inData_25(wire_con_in_stage4[25]), .inData_26(wire_con_in_stage4[26]), .inData_27(wire_con_in_stage4[27]), .inData_28(wire_con_in_stage4[28]), .inData_29(wire_con_in_stage4[29]), .inData_30(wire_con_in_stage4[30]), .inData_31(wire_con_in_stage4[31]), .inData_32(wire_con_in_stage4[32]), .inData_33(wire_con_in_stage4[33]), .inData_34(wire_con_in_stage4[34]), .inData_35(wire_con_in_stage4[35]), .inData_36(wire_con_in_stage4[36]), .inData_37(wire_con_in_stage4[37]), .inData_38(wire_con_in_stage4[38]), .inData_39(wire_con_in_stage4[39]), .inData_40(wire_con_in_stage4[40]), .inData_41(wire_con_in_stage4[41]), .inData_42(wire_con_in_stage4[42]), .inData_43(wire_con_in_stage4[43]), .inData_44(wire_con_in_stage4[44]), .inData_45(wire_con_in_stage4[45]), .inData_46(wire_con_in_stage4[46]), .inData_47(wire_con_in_stage4[47]), .inData_48(wire_con_in_stage4[48]), .inData_49(wire_con_in_stage4[49]), .inData_50(wire_con_in_stage4[50]), .inData_51(wire_con_in_stage4[51]), .inData_52(wire_con_in_stage4[52]), .inData_53(wire_con_in_stage4[53]), .inData_54(wire_con_in_stage4[54]), .inData_55(wire_con_in_stage4[55]), .inData_56(wire_con_in_stage4[56]), .inData_57(wire_con_in_stage4[57]), .inData_58(wire_con_in_stage4[58]), .inData_59(wire_con_in_stage4[59]), .inData_60(wire_con_in_stage4[60]), .inData_61(wire_con_in_stage4[61]), .inData_62(wire_con_in_stage4[62]), .inData_63(wire_con_in_stage4[63]), .inData_64(wire_con_in_stage4[64]), .inData_65(wire_con_in_stage4[65]), .inData_66(wire_con_in_stage4[66]), .inData_67(wire_con_in_stage4[67]), .inData_68(wire_con_in_stage4[68]), .inData_69(wire_con_in_stage4[69]), .inData_70(wire_con_in_stage4[70]), .inData_71(wire_con_in_stage4[71]), .inData_72(wire_con_in_stage4[72]), .inData_73(wire_con_in_stage4[73]), .inData_74(wire_con_in_stage4[74]), .inData_75(wire_con_in_stage4[75]), .inData_76(wire_con_in_stage4[76]), .inData_77(wire_con_in_stage4[77]), .inData_78(wire_con_in_stage4[78]), .inData_79(wire_con_in_stage4[79]), .inData_80(wire_con_in_stage4[80]), .inData_81(wire_con_in_stage4[81]), .inData_82(wire_con_in_stage4[82]), .inData_83(wire_con_in_stage4[83]), .inData_84(wire_con_in_stage4[84]), .inData_85(wire_con_in_stage4[85]), .inData_86(wire_con_in_stage4[86]), .inData_87(wire_con_in_stage4[87]), .inData_88(wire_con_in_stage4[88]), .inData_89(wire_con_in_stage4[89]), .inData_90(wire_con_in_stage4[90]), .inData_91(wire_con_in_stage4[91]), .inData_92(wire_con_in_stage4[92]), .inData_93(wire_con_in_stage4[93]), .inData_94(wire_con_in_stage4[94]), .inData_95(wire_con_in_stage4[95]), .inData_96(wire_con_in_stage4[96]), .inData_97(wire_con_in_stage4[97]), .inData_98(wire_con_in_stage4[98]), .inData_99(wire_con_in_stage4[99]), .inData_100(wire_con_in_stage4[100]), .inData_101(wire_con_in_stage4[101]), .inData_102(wire_con_in_stage4[102]), .inData_103(wire_con_in_stage4[103]), .inData_104(wire_con_in_stage4[104]), .inData_105(wire_con_in_stage4[105]), .inData_106(wire_con_in_stage4[106]), .inData_107(wire_con_in_stage4[107]), .inData_108(wire_con_in_stage4[108]), .inData_109(wire_con_in_stage4[109]), .inData_110(wire_con_in_stage4[110]), .inData_111(wire_con_in_stage4[111]), .inData_112(wire_con_in_stage4[112]), .inData_113(wire_con_in_stage4[113]), .inData_114(wire_con_in_stage4[114]), .inData_115(wire_con_in_stage4[115]), .inData_116(wire_con_in_stage4[116]), .inData_117(wire_con_in_stage4[117]), .inData_118(wire_con_in_stage4[118]), .inData_119(wire_con_in_stage4[119]), .inData_120(wire_con_in_stage4[120]), .inData_121(wire_con_in_stage4[121]), .inData_122(wire_con_in_stage4[122]), .inData_123(wire_con_in_stage4[123]), .inData_124(wire_con_in_stage4[124]), .inData_125(wire_con_in_stage4[125]), .inData_126(wire_con_in_stage4[126]), .inData_127(wire_con_in_stage4[127]), .inData_128(wire_con_in_stage4[128]), .inData_129(wire_con_in_stage4[129]), .inData_130(wire_con_in_stage4[130]), .inData_131(wire_con_in_stage4[131]), .inData_132(wire_con_in_stage4[132]), .inData_133(wire_con_in_stage4[133]), .inData_134(wire_con_in_stage4[134]), .inData_135(wire_con_in_stage4[135]), .inData_136(wire_con_in_stage4[136]), .inData_137(wire_con_in_stage4[137]), .inData_138(wire_con_in_stage4[138]), .inData_139(wire_con_in_stage4[139]), .inData_140(wire_con_in_stage4[140]), .inData_141(wire_con_in_stage4[141]), .inData_142(wire_con_in_stage4[142]), .inData_143(wire_con_in_stage4[143]), .inData_144(wire_con_in_stage4[144]), .inData_145(wire_con_in_stage4[145]), .inData_146(wire_con_in_stage4[146]), .inData_147(wire_con_in_stage4[147]), .inData_148(wire_con_in_stage4[148]), .inData_149(wire_con_in_stage4[149]), .inData_150(wire_con_in_stage4[150]), .inData_151(wire_con_in_stage4[151]), .inData_152(wire_con_in_stage4[152]), .inData_153(wire_con_in_stage4[153]), .inData_154(wire_con_in_stage4[154]), .inData_155(wire_con_in_stage4[155]), .inData_156(wire_con_in_stage4[156]), .inData_157(wire_con_in_stage4[157]), .inData_158(wire_con_in_stage4[158]), .inData_159(wire_con_in_stage4[159]), .inData_160(wire_con_in_stage4[160]), .inData_161(wire_con_in_stage4[161]), .inData_162(wire_con_in_stage4[162]), .inData_163(wire_con_in_stage4[163]), .inData_164(wire_con_in_stage4[164]), .inData_165(wire_con_in_stage4[165]), .inData_166(wire_con_in_stage4[166]), .inData_167(wire_con_in_stage4[167]), .inData_168(wire_con_in_stage4[168]), .inData_169(wire_con_in_stage4[169]), .inData_170(wire_con_in_stage4[170]), .inData_171(wire_con_in_stage4[171]), .inData_172(wire_con_in_stage4[172]), .inData_173(wire_con_in_stage4[173]), .inData_174(wire_con_in_stage4[174]), .inData_175(wire_con_in_stage4[175]), .inData_176(wire_con_in_stage4[176]), .inData_177(wire_con_in_stage4[177]), .inData_178(wire_con_in_stage4[178]), .inData_179(wire_con_in_stage4[179]), .inData_180(wire_con_in_stage4[180]), .inData_181(wire_con_in_stage4[181]), .inData_182(wire_con_in_stage4[182]), .inData_183(wire_con_in_stage4[183]), .inData_184(wire_con_in_stage4[184]), .inData_185(wire_con_in_stage4[185]), .inData_186(wire_con_in_stage4[186]), .inData_187(wire_con_in_stage4[187]), .inData_188(wire_con_in_stage4[188]), .inData_189(wire_con_in_stage4[189]), .inData_190(wire_con_in_stage4[190]), .inData_191(wire_con_in_stage4[191]), .inData_192(wire_con_in_stage4[192]), .inData_193(wire_con_in_stage4[193]), .inData_194(wire_con_in_stage4[194]), .inData_195(wire_con_in_stage4[195]), .inData_196(wire_con_in_stage4[196]), .inData_197(wire_con_in_stage4[197]), .inData_198(wire_con_in_stage4[198]), .inData_199(wire_con_in_stage4[199]), .inData_200(wire_con_in_stage4[200]), .inData_201(wire_con_in_stage4[201]), .inData_202(wire_con_in_stage4[202]), .inData_203(wire_con_in_stage4[203]), .inData_204(wire_con_in_stage4[204]), .inData_205(wire_con_in_stage4[205]), .inData_206(wire_con_in_stage4[206]), .inData_207(wire_con_in_stage4[207]), .inData_208(wire_con_in_stage4[208]), .inData_209(wire_con_in_stage4[209]), .inData_210(wire_con_in_stage4[210]), .inData_211(wire_con_in_stage4[211]), .inData_212(wire_con_in_stage4[212]), .inData_213(wire_con_in_stage4[213]), .inData_214(wire_con_in_stage4[214]), .inData_215(wire_con_in_stage4[215]), .inData_216(wire_con_in_stage4[216]), .inData_217(wire_con_in_stage4[217]), .inData_218(wire_con_in_stage4[218]), .inData_219(wire_con_in_stage4[219]), .inData_220(wire_con_in_stage4[220]), .inData_221(wire_con_in_stage4[221]), .inData_222(wire_con_in_stage4[222]), .inData_223(wire_con_in_stage4[223]), .inData_224(wire_con_in_stage4[224]), .inData_225(wire_con_in_stage4[225]), .inData_226(wire_con_in_stage4[226]), .inData_227(wire_con_in_stage4[227]), .inData_228(wire_con_in_stage4[228]), .inData_229(wire_con_in_stage4[229]), .inData_230(wire_con_in_stage4[230]), .inData_231(wire_con_in_stage4[231]), .inData_232(wire_con_in_stage4[232]), .inData_233(wire_con_in_stage4[233]), .inData_234(wire_con_in_stage4[234]), .inData_235(wire_con_in_stage4[235]), .inData_236(wire_con_in_stage4[236]), .inData_237(wire_con_in_stage4[237]), .inData_238(wire_con_in_stage4[238]), .inData_239(wire_con_in_stage4[239]), .inData_240(wire_con_in_stage4[240]), .inData_241(wire_con_in_stage4[241]), .inData_242(wire_con_in_stage4[242]), .inData_243(wire_con_in_stage4[243]), .inData_244(wire_con_in_stage4[244]), .inData_245(wire_con_in_stage4[245]), .inData_246(wire_con_in_stage4[246]), .inData_247(wire_con_in_stage4[247]), .inData_248(wire_con_in_stage4[248]), .inData_249(wire_con_in_stage4[249]), .inData_250(wire_con_in_stage4[250]), .inData_251(wire_con_in_stage4[251]), .inData_252(wire_con_in_stage4[252]), .inData_253(wire_con_in_stage4[253]), .inData_254(wire_con_in_stage4[254]), .inData_255(wire_con_in_stage4[255]), 
        .outData_0(wire_con_out_stage4[0]), .outData_1(wire_con_out_stage4[1]), .outData_2(wire_con_out_stage4[2]), .outData_3(wire_con_out_stage4[3]), .outData_4(wire_con_out_stage4[4]), .outData_5(wire_con_out_stage4[5]), .outData_6(wire_con_out_stage4[6]), .outData_7(wire_con_out_stage4[7]), .outData_8(wire_con_out_stage4[8]), .outData_9(wire_con_out_stage4[9]), .outData_10(wire_con_out_stage4[10]), .outData_11(wire_con_out_stage4[11]), .outData_12(wire_con_out_stage4[12]), .outData_13(wire_con_out_stage4[13]), .outData_14(wire_con_out_stage4[14]), .outData_15(wire_con_out_stage4[15]), .outData_16(wire_con_out_stage4[16]), .outData_17(wire_con_out_stage4[17]), .outData_18(wire_con_out_stage4[18]), .outData_19(wire_con_out_stage4[19]), .outData_20(wire_con_out_stage4[20]), .outData_21(wire_con_out_stage4[21]), .outData_22(wire_con_out_stage4[22]), .outData_23(wire_con_out_stage4[23]), .outData_24(wire_con_out_stage4[24]), .outData_25(wire_con_out_stage4[25]), .outData_26(wire_con_out_stage4[26]), .outData_27(wire_con_out_stage4[27]), .outData_28(wire_con_out_stage4[28]), .outData_29(wire_con_out_stage4[29]), .outData_30(wire_con_out_stage4[30]), .outData_31(wire_con_out_stage4[31]), .outData_32(wire_con_out_stage4[32]), .outData_33(wire_con_out_stage4[33]), .outData_34(wire_con_out_stage4[34]), .outData_35(wire_con_out_stage4[35]), .outData_36(wire_con_out_stage4[36]), .outData_37(wire_con_out_stage4[37]), .outData_38(wire_con_out_stage4[38]), .outData_39(wire_con_out_stage4[39]), .outData_40(wire_con_out_stage4[40]), .outData_41(wire_con_out_stage4[41]), .outData_42(wire_con_out_stage4[42]), .outData_43(wire_con_out_stage4[43]), .outData_44(wire_con_out_stage4[44]), .outData_45(wire_con_out_stage4[45]), .outData_46(wire_con_out_stage4[46]), .outData_47(wire_con_out_stage4[47]), .outData_48(wire_con_out_stage4[48]), .outData_49(wire_con_out_stage4[49]), .outData_50(wire_con_out_stage4[50]), .outData_51(wire_con_out_stage4[51]), .outData_52(wire_con_out_stage4[52]), .outData_53(wire_con_out_stage4[53]), .outData_54(wire_con_out_stage4[54]), .outData_55(wire_con_out_stage4[55]), .outData_56(wire_con_out_stage4[56]), .outData_57(wire_con_out_stage4[57]), .outData_58(wire_con_out_stage4[58]), .outData_59(wire_con_out_stage4[59]), .outData_60(wire_con_out_stage4[60]), .outData_61(wire_con_out_stage4[61]), .outData_62(wire_con_out_stage4[62]), .outData_63(wire_con_out_stage4[63]), .outData_64(wire_con_out_stage4[64]), .outData_65(wire_con_out_stage4[65]), .outData_66(wire_con_out_stage4[66]), .outData_67(wire_con_out_stage4[67]), .outData_68(wire_con_out_stage4[68]), .outData_69(wire_con_out_stage4[69]), .outData_70(wire_con_out_stage4[70]), .outData_71(wire_con_out_stage4[71]), .outData_72(wire_con_out_stage4[72]), .outData_73(wire_con_out_stage4[73]), .outData_74(wire_con_out_stage4[74]), .outData_75(wire_con_out_stage4[75]), .outData_76(wire_con_out_stage4[76]), .outData_77(wire_con_out_stage4[77]), .outData_78(wire_con_out_stage4[78]), .outData_79(wire_con_out_stage4[79]), .outData_80(wire_con_out_stage4[80]), .outData_81(wire_con_out_stage4[81]), .outData_82(wire_con_out_stage4[82]), .outData_83(wire_con_out_stage4[83]), .outData_84(wire_con_out_stage4[84]), .outData_85(wire_con_out_stage4[85]), .outData_86(wire_con_out_stage4[86]), .outData_87(wire_con_out_stage4[87]), .outData_88(wire_con_out_stage4[88]), .outData_89(wire_con_out_stage4[89]), .outData_90(wire_con_out_stage4[90]), .outData_91(wire_con_out_stage4[91]), .outData_92(wire_con_out_stage4[92]), .outData_93(wire_con_out_stage4[93]), .outData_94(wire_con_out_stage4[94]), .outData_95(wire_con_out_stage4[95]), .outData_96(wire_con_out_stage4[96]), .outData_97(wire_con_out_stage4[97]), .outData_98(wire_con_out_stage4[98]), .outData_99(wire_con_out_stage4[99]), .outData_100(wire_con_out_stage4[100]), .outData_101(wire_con_out_stage4[101]), .outData_102(wire_con_out_stage4[102]), .outData_103(wire_con_out_stage4[103]), .outData_104(wire_con_out_stage4[104]), .outData_105(wire_con_out_stage4[105]), .outData_106(wire_con_out_stage4[106]), .outData_107(wire_con_out_stage4[107]), .outData_108(wire_con_out_stage4[108]), .outData_109(wire_con_out_stage4[109]), .outData_110(wire_con_out_stage4[110]), .outData_111(wire_con_out_stage4[111]), .outData_112(wire_con_out_stage4[112]), .outData_113(wire_con_out_stage4[113]), .outData_114(wire_con_out_stage4[114]), .outData_115(wire_con_out_stage4[115]), .outData_116(wire_con_out_stage4[116]), .outData_117(wire_con_out_stage4[117]), .outData_118(wire_con_out_stage4[118]), .outData_119(wire_con_out_stage4[119]), .outData_120(wire_con_out_stage4[120]), .outData_121(wire_con_out_stage4[121]), .outData_122(wire_con_out_stage4[122]), .outData_123(wire_con_out_stage4[123]), .outData_124(wire_con_out_stage4[124]), .outData_125(wire_con_out_stage4[125]), .outData_126(wire_con_out_stage4[126]), .outData_127(wire_con_out_stage4[127]), .outData_128(wire_con_out_stage4[128]), .outData_129(wire_con_out_stage4[129]), .outData_130(wire_con_out_stage4[130]), .outData_131(wire_con_out_stage4[131]), .outData_132(wire_con_out_stage4[132]), .outData_133(wire_con_out_stage4[133]), .outData_134(wire_con_out_stage4[134]), .outData_135(wire_con_out_stage4[135]), .outData_136(wire_con_out_stage4[136]), .outData_137(wire_con_out_stage4[137]), .outData_138(wire_con_out_stage4[138]), .outData_139(wire_con_out_stage4[139]), .outData_140(wire_con_out_stage4[140]), .outData_141(wire_con_out_stage4[141]), .outData_142(wire_con_out_stage4[142]), .outData_143(wire_con_out_stage4[143]), .outData_144(wire_con_out_stage4[144]), .outData_145(wire_con_out_stage4[145]), .outData_146(wire_con_out_stage4[146]), .outData_147(wire_con_out_stage4[147]), .outData_148(wire_con_out_stage4[148]), .outData_149(wire_con_out_stage4[149]), .outData_150(wire_con_out_stage4[150]), .outData_151(wire_con_out_stage4[151]), .outData_152(wire_con_out_stage4[152]), .outData_153(wire_con_out_stage4[153]), .outData_154(wire_con_out_stage4[154]), .outData_155(wire_con_out_stage4[155]), .outData_156(wire_con_out_stage4[156]), .outData_157(wire_con_out_stage4[157]), .outData_158(wire_con_out_stage4[158]), .outData_159(wire_con_out_stage4[159]), .outData_160(wire_con_out_stage4[160]), .outData_161(wire_con_out_stage4[161]), .outData_162(wire_con_out_stage4[162]), .outData_163(wire_con_out_stage4[163]), .outData_164(wire_con_out_stage4[164]), .outData_165(wire_con_out_stage4[165]), .outData_166(wire_con_out_stage4[166]), .outData_167(wire_con_out_stage4[167]), .outData_168(wire_con_out_stage4[168]), .outData_169(wire_con_out_stage4[169]), .outData_170(wire_con_out_stage4[170]), .outData_171(wire_con_out_stage4[171]), .outData_172(wire_con_out_stage4[172]), .outData_173(wire_con_out_stage4[173]), .outData_174(wire_con_out_stage4[174]), .outData_175(wire_con_out_stage4[175]), .outData_176(wire_con_out_stage4[176]), .outData_177(wire_con_out_stage4[177]), .outData_178(wire_con_out_stage4[178]), .outData_179(wire_con_out_stage4[179]), .outData_180(wire_con_out_stage4[180]), .outData_181(wire_con_out_stage4[181]), .outData_182(wire_con_out_stage4[182]), .outData_183(wire_con_out_stage4[183]), .outData_184(wire_con_out_stage4[184]), .outData_185(wire_con_out_stage4[185]), .outData_186(wire_con_out_stage4[186]), .outData_187(wire_con_out_stage4[187]), .outData_188(wire_con_out_stage4[188]), .outData_189(wire_con_out_stage4[189]), .outData_190(wire_con_out_stage4[190]), .outData_191(wire_con_out_stage4[191]), .outData_192(wire_con_out_stage4[192]), .outData_193(wire_con_out_stage4[193]), .outData_194(wire_con_out_stage4[194]), .outData_195(wire_con_out_stage4[195]), .outData_196(wire_con_out_stage4[196]), .outData_197(wire_con_out_stage4[197]), .outData_198(wire_con_out_stage4[198]), .outData_199(wire_con_out_stage4[199]), .outData_200(wire_con_out_stage4[200]), .outData_201(wire_con_out_stage4[201]), .outData_202(wire_con_out_stage4[202]), .outData_203(wire_con_out_stage4[203]), .outData_204(wire_con_out_stage4[204]), .outData_205(wire_con_out_stage4[205]), .outData_206(wire_con_out_stage4[206]), .outData_207(wire_con_out_stage4[207]), .outData_208(wire_con_out_stage4[208]), .outData_209(wire_con_out_stage4[209]), .outData_210(wire_con_out_stage4[210]), .outData_211(wire_con_out_stage4[211]), .outData_212(wire_con_out_stage4[212]), .outData_213(wire_con_out_stage4[213]), .outData_214(wire_con_out_stage4[214]), .outData_215(wire_con_out_stage4[215]), .outData_216(wire_con_out_stage4[216]), .outData_217(wire_con_out_stage4[217]), .outData_218(wire_con_out_stage4[218]), .outData_219(wire_con_out_stage4[219]), .outData_220(wire_con_out_stage4[220]), .outData_221(wire_con_out_stage4[221]), .outData_222(wire_con_out_stage4[222]), .outData_223(wire_con_out_stage4[223]), .outData_224(wire_con_out_stage4[224]), .outData_225(wire_con_out_stage4[225]), .outData_226(wire_con_out_stage4[226]), .outData_227(wire_con_out_stage4[227]), .outData_228(wire_con_out_stage4[228]), .outData_229(wire_con_out_stage4[229]), .outData_230(wire_con_out_stage4[230]), .outData_231(wire_con_out_stage4[231]), .outData_232(wire_con_out_stage4[232]), .outData_233(wire_con_out_stage4[233]), .outData_234(wire_con_out_stage4[234]), .outData_235(wire_con_out_stage4[235]), .outData_236(wire_con_out_stage4[236]), .outData_237(wire_con_out_stage4[237]), .outData_238(wire_con_out_stage4[238]), .outData_239(wire_con_out_stage4[239]), .outData_240(wire_con_out_stage4[240]), .outData_241(wire_con_out_stage4[241]), .outData_242(wire_con_out_stage4[242]), .outData_243(wire_con_out_stage4[243]), .outData_244(wire_con_out_stage4[244]), .outData_245(wire_con_out_stage4[245]), .outData_246(wire_con_out_stage4[246]), .outData_247(wire_con_out_stage4[247]), .outData_248(wire_con_out_stage4[248]), .outData_249(wire_con_out_stage4[249]), .outData_250(wire_con_out_stage4[250]), .outData_251(wire_con_out_stage4[251]), .outData_252(wire_con_out_stage4[252]), .outData_253(wire_con_out_stage4[253]), .outData_254(wire_con_out_stage4[254]), .outData_255(wire_con_out_stage4[255]), 
        .in_start(con_in_start_stage4), .out_start(in_start_stage5), .clk(clk), .rst(rst)); 

  
  assign wire_ctrl_stage4[0] = counter_w[3]; 
  assign wire_ctrl_stage4[1] = counter_w[3]; 
  assign wire_ctrl_stage4[2] = counter_w[3]; 
  assign wire_ctrl_stage4[3] = counter_w[3]; 
  assign wire_ctrl_stage4[4] = counter_w[3]; 
  assign wire_ctrl_stage4[5] = counter_w[3]; 
  assign wire_ctrl_stage4[6] = counter_w[3]; 
  assign wire_ctrl_stage4[7] = counter_w[3]; 
  assign wire_ctrl_stage4[8] = counter_w[3]; 
  assign wire_ctrl_stage4[9] = counter_w[3]; 
  assign wire_ctrl_stage4[10] = counter_w[3]; 
  assign wire_ctrl_stage4[11] = counter_w[3]; 
  assign wire_ctrl_stage4[12] = counter_w[3]; 
  assign wire_ctrl_stage4[13] = counter_w[3]; 
  assign wire_ctrl_stage4[14] = counter_w[3]; 
  assign wire_ctrl_stage4[15] = counter_w[3]; 
  assign wire_ctrl_stage4[16] = counter_w[3]; 
  assign wire_ctrl_stage4[17] = counter_w[3]; 
  assign wire_ctrl_stage4[18] = counter_w[3]; 
  assign wire_ctrl_stage4[19] = counter_w[3]; 
  assign wire_ctrl_stage4[20] = counter_w[3]; 
  assign wire_ctrl_stage4[21] = counter_w[3]; 
  assign wire_ctrl_stage4[22] = counter_w[3]; 
  assign wire_ctrl_stage4[23] = counter_w[3]; 
  assign wire_ctrl_stage4[24] = counter_w[3]; 
  assign wire_ctrl_stage4[25] = counter_w[3]; 
  assign wire_ctrl_stage4[26] = counter_w[3]; 
  assign wire_ctrl_stage4[27] = counter_w[3]; 
  assign wire_ctrl_stage4[28] = counter_w[3]; 
  assign wire_ctrl_stage4[29] = counter_w[3]; 
  assign wire_ctrl_stage4[30] = counter_w[3]; 
  assign wire_ctrl_stage4[31] = counter_w[3]; 
  assign wire_ctrl_stage4[32] = counter_w[3]; 
  assign wire_ctrl_stage4[33] = counter_w[3]; 
  assign wire_ctrl_stage4[34] = counter_w[3]; 
  assign wire_ctrl_stage4[35] = counter_w[3]; 
  assign wire_ctrl_stage4[36] = counter_w[3]; 
  assign wire_ctrl_stage4[37] = counter_w[3]; 
  assign wire_ctrl_stage4[38] = counter_w[3]; 
  assign wire_ctrl_stage4[39] = counter_w[3]; 
  assign wire_ctrl_stage4[40] = counter_w[3]; 
  assign wire_ctrl_stage4[41] = counter_w[3]; 
  assign wire_ctrl_stage4[42] = counter_w[3]; 
  assign wire_ctrl_stage4[43] = counter_w[3]; 
  assign wire_ctrl_stage4[44] = counter_w[3]; 
  assign wire_ctrl_stage4[45] = counter_w[3]; 
  assign wire_ctrl_stage4[46] = counter_w[3]; 
  assign wire_ctrl_stage4[47] = counter_w[3]; 
  assign wire_ctrl_stage4[48] = counter_w[3]; 
  assign wire_ctrl_stage4[49] = counter_w[3]; 
  assign wire_ctrl_stage4[50] = counter_w[3]; 
  assign wire_ctrl_stage4[51] = counter_w[3]; 
  assign wire_ctrl_stage4[52] = counter_w[3]; 
  assign wire_ctrl_stage4[53] = counter_w[3]; 
  assign wire_ctrl_stage4[54] = counter_w[3]; 
  assign wire_ctrl_stage4[55] = counter_w[3]; 
  assign wire_ctrl_stage4[56] = counter_w[3]; 
  assign wire_ctrl_stage4[57] = counter_w[3]; 
  assign wire_ctrl_stage4[58] = counter_w[3]; 
  assign wire_ctrl_stage4[59] = counter_w[3]; 
  assign wire_ctrl_stage4[60] = counter_w[3]; 
  assign wire_ctrl_stage4[61] = counter_w[3]; 
  assign wire_ctrl_stage4[62] = counter_w[3]; 
  assign wire_ctrl_stage4[63] = counter_w[3]; 
  assign wire_ctrl_stage4[64] = counter_w[3]; 
  assign wire_ctrl_stage4[65] = counter_w[3]; 
  assign wire_ctrl_stage4[66] = counter_w[3]; 
  assign wire_ctrl_stage4[67] = counter_w[3]; 
  assign wire_ctrl_stage4[68] = counter_w[3]; 
  assign wire_ctrl_stage4[69] = counter_w[3]; 
  assign wire_ctrl_stage4[70] = counter_w[3]; 
  assign wire_ctrl_stage4[71] = counter_w[3]; 
  assign wire_ctrl_stage4[72] = counter_w[3]; 
  assign wire_ctrl_stage4[73] = counter_w[3]; 
  assign wire_ctrl_stage4[74] = counter_w[3]; 
  assign wire_ctrl_stage4[75] = counter_w[3]; 
  assign wire_ctrl_stage4[76] = counter_w[3]; 
  assign wire_ctrl_stage4[77] = counter_w[3]; 
  assign wire_ctrl_stage4[78] = counter_w[3]; 
  assign wire_ctrl_stage4[79] = counter_w[3]; 
  assign wire_ctrl_stage4[80] = counter_w[3]; 
  assign wire_ctrl_stage4[81] = counter_w[3]; 
  assign wire_ctrl_stage4[82] = counter_w[3]; 
  assign wire_ctrl_stage4[83] = counter_w[3]; 
  assign wire_ctrl_stage4[84] = counter_w[3]; 
  assign wire_ctrl_stage4[85] = counter_w[3]; 
  assign wire_ctrl_stage4[86] = counter_w[3]; 
  assign wire_ctrl_stage4[87] = counter_w[3]; 
  assign wire_ctrl_stage4[88] = counter_w[3]; 
  assign wire_ctrl_stage4[89] = counter_w[3]; 
  assign wire_ctrl_stage4[90] = counter_w[3]; 
  assign wire_ctrl_stage4[91] = counter_w[3]; 
  assign wire_ctrl_stage4[92] = counter_w[3]; 
  assign wire_ctrl_stage4[93] = counter_w[3]; 
  assign wire_ctrl_stage4[94] = counter_w[3]; 
  assign wire_ctrl_stage4[95] = counter_w[3]; 
  assign wire_ctrl_stage4[96] = counter_w[3]; 
  assign wire_ctrl_stage4[97] = counter_w[3]; 
  assign wire_ctrl_stage4[98] = counter_w[3]; 
  assign wire_ctrl_stage4[99] = counter_w[3]; 
  assign wire_ctrl_stage4[100] = counter_w[3]; 
  assign wire_ctrl_stage4[101] = counter_w[3]; 
  assign wire_ctrl_stage4[102] = counter_w[3]; 
  assign wire_ctrl_stage4[103] = counter_w[3]; 
  assign wire_ctrl_stage4[104] = counter_w[3]; 
  assign wire_ctrl_stage4[105] = counter_w[3]; 
  assign wire_ctrl_stage4[106] = counter_w[3]; 
  assign wire_ctrl_stage4[107] = counter_w[3]; 
  assign wire_ctrl_stage4[108] = counter_w[3]; 
  assign wire_ctrl_stage4[109] = counter_w[3]; 
  assign wire_ctrl_stage4[110] = counter_w[3]; 
  assign wire_ctrl_stage4[111] = counter_w[3]; 
  assign wire_ctrl_stage4[112] = counter_w[3]; 
  assign wire_ctrl_stage4[113] = counter_w[3]; 
  assign wire_ctrl_stage4[114] = counter_w[3]; 
  assign wire_ctrl_stage4[115] = counter_w[3]; 
  assign wire_ctrl_stage4[116] = counter_w[3]; 
  assign wire_ctrl_stage4[117] = counter_w[3]; 
  assign wire_ctrl_stage4[118] = counter_w[3]; 
  assign wire_ctrl_stage4[119] = counter_w[3]; 
  assign wire_ctrl_stage4[120] = counter_w[3]; 
  assign wire_ctrl_stage4[121] = counter_w[3]; 
  assign wire_ctrl_stage4[122] = counter_w[3]; 
  assign wire_ctrl_stage4[123] = counter_w[3]; 
  assign wire_ctrl_stage4[124] = counter_w[3]; 
  assign wire_ctrl_stage4[125] = counter_w[3]; 
  assign wire_ctrl_stage4[126] = counter_w[3]; 
  assign wire_ctrl_stage4[127] = counter_w[3]; 
  wire [DATA_WIDTH-1:0] wire_con_in_stage5[255:0];
  wire [DATA_WIDTH-1:0] wire_con_out_stage5[255:0];
  wire [127:0] wire_ctrl_stage5;

  switches_stage_st5_0_L switch_stage_5(
        .inData_0(wire_con_out_stage4[0]), .inData_1(wire_con_out_stage4[1]), .inData_2(wire_con_out_stage4[2]), .inData_3(wire_con_out_stage4[3]), .inData_4(wire_con_out_stage4[4]), .inData_5(wire_con_out_stage4[5]), .inData_6(wire_con_out_stage4[6]), .inData_7(wire_con_out_stage4[7]), .inData_8(wire_con_out_stage4[8]), .inData_9(wire_con_out_stage4[9]), .inData_10(wire_con_out_stage4[10]), .inData_11(wire_con_out_stage4[11]), .inData_12(wire_con_out_stage4[12]), .inData_13(wire_con_out_stage4[13]), .inData_14(wire_con_out_stage4[14]), .inData_15(wire_con_out_stage4[15]), .inData_16(wire_con_out_stage4[16]), .inData_17(wire_con_out_stage4[17]), .inData_18(wire_con_out_stage4[18]), .inData_19(wire_con_out_stage4[19]), .inData_20(wire_con_out_stage4[20]), .inData_21(wire_con_out_stage4[21]), .inData_22(wire_con_out_stage4[22]), .inData_23(wire_con_out_stage4[23]), .inData_24(wire_con_out_stage4[24]), .inData_25(wire_con_out_stage4[25]), .inData_26(wire_con_out_stage4[26]), .inData_27(wire_con_out_stage4[27]), .inData_28(wire_con_out_stage4[28]), .inData_29(wire_con_out_stage4[29]), .inData_30(wire_con_out_stage4[30]), .inData_31(wire_con_out_stage4[31]), .inData_32(wire_con_out_stage4[32]), .inData_33(wire_con_out_stage4[33]), .inData_34(wire_con_out_stage4[34]), .inData_35(wire_con_out_stage4[35]), .inData_36(wire_con_out_stage4[36]), .inData_37(wire_con_out_stage4[37]), .inData_38(wire_con_out_stage4[38]), .inData_39(wire_con_out_stage4[39]), .inData_40(wire_con_out_stage4[40]), .inData_41(wire_con_out_stage4[41]), .inData_42(wire_con_out_stage4[42]), .inData_43(wire_con_out_stage4[43]), .inData_44(wire_con_out_stage4[44]), .inData_45(wire_con_out_stage4[45]), .inData_46(wire_con_out_stage4[46]), .inData_47(wire_con_out_stage4[47]), .inData_48(wire_con_out_stage4[48]), .inData_49(wire_con_out_stage4[49]), .inData_50(wire_con_out_stage4[50]), .inData_51(wire_con_out_stage4[51]), .inData_52(wire_con_out_stage4[52]), .inData_53(wire_con_out_stage4[53]), .inData_54(wire_con_out_stage4[54]), .inData_55(wire_con_out_stage4[55]), .inData_56(wire_con_out_stage4[56]), .inData_57(wire_con_out_stage4[57]), .inData_58(wire_con_out_stage4[58]), .inData_59(wire_con_out_stage4[59]), .inData_60(wire_con_out_stage4[60]), .inData_61(wire_con_out_stage4[61]), .inData_62(wire_con_out_stage4[62]), .inData_63(wire_con_out_stage4[63]), .inData_64(wire_con_out_stage4[64]), .inData_65(wire_con_out_stage4[65]), .inData_66(wire_con_out_stage4[66]), .inData_67(wire_con_out_stage4[67]), .inData_68(wire_con_out_stage4[68]), .inData_69(wire_con_out_stage4[69]), .inData_70(wire_con_out_stage4[70]), .inData_71(wire_con_out_stage4[71]), .inData_72(wire_con_out_stage4[72]), .inData_73(wire_con_out_stage4[73]), .inData_74(wire_con_out_stage4[74]), .inData_75(wire_con_out_stage4[75]), .inData_76(wire_con_out_stage4[76]), .inData_77(wire_con_out_stage4[77]), .inData_78(wire_con_out_stage4[78]), .inData_79(wire_con_out_stage4[79]), .inData_80(wire_con_out_stage4[80]), .inData_81(wire_con_out_stage4[81]), .inData_82(wire_con_out_stage4[82]), .inData_83(wire_con_out_stage4[83]), .inData_84(wire_con_out_stage4[84]), .inData_85(wire_con_out_stage4[85]), .inData_86(wire_con_out_stage4[86]), .inData_87(wire_con_out_stage4[87]), .inData_88(wire_con_out_stage4[88]), .inData_89(wire_con_out_stage4[89]), .inData_90(wire_con_out_stage4[90]), .inData_91(wire_con_out_stage4[91]), .inData_92(wire_con_out_stage4[92]), .inData_93(wire_con_out_stage4[93]), .inData_94(wire_con_out_stage4[94]), .inData_95(wire_con_out_stage4[95]), .inData_96(wire_con_out_stage4[96]), .inData_97(wire_con_out_stage4[97]), .inData_98(wire_con_out_stage4[98]), .inData_99(wire_con_out_stage4[99]), .inData_100(wire_con_out_stage4[100]), .inData_101(wire_con_out_stage4[101]), .inData_102(wire_con_out_stage4[102]), .inData_103(wire_con_out_stage4[103]), .inData_104(wire_con_out_stage4[104]), .inData_105(wire_con_out_stage4[105]), .inData_106(wire_con_out_stage4[106]), .inData_107(wire_con_out_stage4[107]), .inData_108(wire_con_out_stage4[108]), .inData_109(wire_con_out_stage4[109]), .inData_110(wire_con_out_stage4[110]), .inData_111(wire_con_out_stage4[111]), .inData_112(wire_con_out_stage4[112]), .inData_113(wire_con_out_stage4[113]), .inData_114(wire_con_out_stage4[114]), .inData_115(wire_con_out_stage4[115]), .inData_116(wire_con_out_stage4[116]), .inData_117(wire_con_out_stage4[117]), .inData_118(wire_con_out_stage4[118]), .inData_119(wire_con_out_stage4[119]), .inData_120(wire_con_out_stage4[120]), .inData_121(wire_con_out_stage4[121]), .inData_122(wire_con_out_stage4[122]), .inData_123(wire_con_out_stage4[123]), .inData_124(wire_con_out_stage4[124]), .inData_125(wire_con_out_stage4[125]), .inData_126(wire_con_out_stage4[126]), .inData_127(wire_con_out_stage4[127]), .inData_128(wire_con_out_stage4[128]), .inData_129(wire_con_out_stage4[129]), .inData_130(wire_con_out_stage4[130]), .inData_131(wire_con_out_stage4[131]), .inData_132(wire_con_out_stage4[132]), .inData_133(wire_con_out_stage4[133]), .inData_134(wire_con_out_stage4[134]), .inData_135(wire_con_out_stage4[135]), .inData_136(wire_con_out_stage4[136]), .inData_137(wire_con_out_stage4[137]), .inData_138(wire_con_out_stage4[138]), .inData_139(wire_con_out_stage4[139]), .inData_140(wire_con_out_stage4[140]), .inData_141(wire_con_out_stage4[141]), .inData_142(wire_con_out_stage4[142]), .inData_143(wire_con_out_stage4[143]), .inData_144(wire_con_out_stage4[144]), .inData_145(wire_con_out_stage4[145]), .inData_146(wire_con_out_stage4[146]), .inData_147(wire_con_out_stage4[147]), .inData_148(wire_con_out_stage4[148]), .inData_149(wire_con_out_stage4[149]), .inData_150(wire_con_out_stage4[150]), .inData_151(wire_con_out_stage4[151]), .inData_152(wire_con_out_stage4[152]), .inData_153(wire_con_out_stage4[153]), .inData_154(wire_con_out_stage4[154]), .inData_155(wire_con_out_stage4[155]), .inData_156(wire_con_out_stage4[156]), .inData_157(wire_con_out_stage4[157]), .inData_158(wire_con_out_stage4[158]), .inData_159(wire_con_out_stage4[159]), .inData_160(wire_con_out_stage4[160]), .inData_161(wire_con_out_stage4[161]), .inData_162(wire_con_out_stage4[162]), .inData_163(wire_con_out_stage4[163]), .inData_164(wire_con_out_stage4[164]), .inData_165(wire_con_out_stage4[165]), .inData_166(wire_con_out_stage4[166]), .inData_167(wire_con_out_stage4[167]), .inData_168(wire_con_out_stage4[168]), .inData_169(wire_con_out_stage4[169]), .inData_170(wire_con_out_stage4[170]), .inData_171(wire_con_out_stage4[171]), .inData_172(wire_con_out_stage4[172]), .inData_173(wire_con_out_stage4[173]), .inData_174(wire_con_out_stage4[174]), .inData_175(wire_con_out_stage4[175]), .inData_176(wire_con_out_stage4[176]), .inData_177(wire_con_out_stage4[177]), .inData_178(wire_con_out_stage4[178]), .inData_179(wire_con_out_stage4[179]), .inData_180(wire_con_out_stage4[180]), .inData_181(wire_con_out_stage4[181]), .inData_182(wire_con_out_stage4[182]), .inData_183(wire_con_out_stage4[183]), .inData_184(wire_con_out_stage4[184]), .inData_185(wire_con_out_stage4[185]), .inData_186(wire_con_out_stage4[186]), .inData_187(wire_con_out_stage4[187]), .inData_188(wire_con_out_stage4[188]), .inData_189(wire_con_out_stage4[189]), .inData_190(wire_con_out_stage4[190]), .inData_191(wire_con_out_stage4[191]), .inData_192(wire_con_out_stage4[192]), .inData_193(wire_con_out_stage4[193]), .inData_194(wire_con_out_stage4[194]), .inData_195(wire_con_out_stage4[195]), .inData_196(wire_con_out_stage4[196]), .inData_197(wire_con_out_stage4[197]), .inData_198(wire_con_out_stage4[198]), .inData_199(wire_con_out_stage4[199]), .inData_200(wire_con_out_stage4[200]), .inData_201(wire_con_out_stage4[201]), .inData_202(wire_con_out_stage4[202]), .inData_203(wire_con_out_stage4[203]), .inData_204(wire_con_out_stage4[204]), .inData_205(wire_con_out_stage4[205]), .inData_206(wire_con_out_stage4[206]), .inData_207(wire_con_out_stage4[207]), .inData_208(wire_con_out_stage4[208]), .inData_209(wire_con_out_stage4[209]), .inData_210(wire_con_out_stage4[210]), .inData_211(wire_con_out_stage4[211]), .inData_212(wire_con_out_stage4[212]), .inData_213(wire_con_out_stage4[213]), .inData_214(wire_con_out_stage4[214]), .inData_215(wire_con_out_stage4[215]), .inData_216(wire_con_out_stage4[216]), .inData_217(wire_con_out_stage4[217]), .inData_218(wire_con_out_stage4[218]), .inData_219(wire_con_out_stage4[219]), .inData_220(wire_con_out_stage4[220]), .inData_221(wire_con_out_stage4[221]), .inData_222(wire_con_out_stage4[222]), .inData_223(wire_con_out_stage4[223]), .inData_224(wire_con_out_stage4[224]), .inData_225(wire_con_out_stage4[225]), .inData_226(wire_con_out_stage4[226]), .inData_227(wire_con_out_stage4[227]), .inData_228(wire_con_out_stage4[228]), .inData_229(wire_con_out_stage4[229]), .inData_230(wire_con_out_stage4[230]), .inData_231(wire_con_out_stage4[231]), .inData_232(wire_con_out_stage4[232]), .inData_233(wire_con_out_stage4[233]), .inData_234(wire_con_out_stage4[234]), .inData_235(wire_con_out_stage4[235]), .inData_236(wire_con_out_stage4[236]), .inData_237(wire_con_out_stage4[237]), .inData_238(wire_con_out_stage4[238]), .inData_239(wire_con_out_stage4[239]), .inData_240(wire_con_out_stage4[240]), .inData_241(wire_con_out_stage4[241]), .inData_242(wire_con_out_stage4[242]), .inData_243(wire_con_out_stage4[243]), .inData_244(wire_con_out_stage4[244]), .inData_245(wire_con_out_stage4[245]), .inData_246(wire_con_out_stage4[246]), .inData_247(wire_con_out_stage4[247]), .inData_248(wire_con_out_stage4[248]), .inData_249(wire_con_out_stage4[249]), .inData_250(wire_con_out_stage4[250]), .inData_251(wire_con_out_stage4[251]), .inData_252(wire_con_out_stage4[252]), .inData_253(wire_con_out_stage4[253]), .inData_254(wire_con_out_stage4[254]), .inData_255(wire_con_out_stage4[255]), 
        .outData_0(wire_con_in_stage5[0]), .outData_1(wire_con_in_stage5[1]), .outData_2(wire_con_in_stage5[2]), .outData_3(wire_con_in_stage5[3]), .outData_4(wire_con_in_stage5[4]), .outData_5(wire_con_in_stage5[5]), .outData_6(wire_con_in_stage5[6]), .outData_7(wire_con_in_stage5[7]), .outData_8(wire_con_in_stage5[8]), .outData_9(wire_con_in_stage5[9]), .outData_10(wire_con_in_stage5[10]), .outData_11(wire_con_in_stage5[11]), .outData_12(wire_con_in_stage5[12]), .outData_13(wire_con_in_stage5[13]), .outData_14(wire_con_in_stage5[14]), .outData_15(wire_con_in_stage5[15]), .outData_16(wire_con_in_stage5[16]), .outData_17(wire_con_in_stage5[17]), .outData_18(wire_con_in_stage5[18]), .outData_19(wire_con_in_stage5[19]), .outData_20(wire_con_in_stage5[20]), .outData_21(wire_con_in_stage5[21]), .outData_22(wire_con_in_stage5[22]), .outData_23(wire_con_in_stage5[23]), .outData_24(wire_con_in_stage5[24]), .outData_25(wire_con_in_stage5[25]), .outData_26(wire_con_in_stage5[26]), .outData_27(wire_con_in_stage5[27]), .outData_28(wire_con_in_stage5[28]), .outData_29(wire_con_in_stage5[29]), .outData_30(wire_con_in_stage5[30]), .outData_31(wire_con_in_stage5[31]), .outData_32(wire_con_in_stage5[32]), .outData_33(wire_con_in_stage5[33]), .outData_34(wire_con_in_stage5[34]), .outData_35(wire_con_in_stage5[35]), .outData_36(wire_con_in_stage5[36]), .outData_37(wire_con_in_stage5[37]), .outData_38(wire_con_in_stage5[38]), .outData_39(wire_con_in_stage5[39]), .outData_40(wire_con_in_stage5[40]), .outData_41(wire_con_in_stage5[41]), .outData_42(wire_con_in_stage5[42]), .outData_43(wire_con_in_stage5[43]), .outData_44(wire_con_in_stage5[44]), .outData_45(wire_con_in_stage5[45]), .outData_46(wire_con_in_stage5[46]), .outData_47(wire_con_in_stage5[47]), .outData_48(wire_con_in_stage5[48]), .outData_49(wire_con_in_stage5[49]), .outData_50(wire_con_in_stage5[50]), .outData_51(wire_con_in_stage5[51]), .outData_52(wire_con_in_stage5[52]), .outData_53(wire_con_in_stage5[53]), .outData_54(wire_con_in_stage5[54]), .outData_55(wire_con_in_stage5[55]), .outData_56(wire_con_in_stage5[56]), .outData_57(wire_con_in_stage5[57]), .outData_58(wire_con_in_stage5[58]), .outData_59(wire_con_in_stage5[59]), .outData_60(wire_con_in_stage5[60]), .outData_61(wire_con_in_stage5[61]), .outData_62(wire_con_in_stage5[62]), .outData_63(wire_con_in_stage5[63]), .outData_64(wire_con_in_stage5[64]), .outData_65(wire_con_in_stage5[65]), .outData_66(wire_con_in_stage5[66]), .outData_67(wire_con_in_stage5[67]), .outData_68(wire_con_in_stage5[68]), .outData_69(wire_con_in_stage5[69]), .outData_70(wire_con_in_stage5[70]), .outData_71(wire_con_in_stage5[71]), .outData_72(wire_con_in_stage5[72]), .outData_73(wire_con_in_stage5[73]), .outData_74(wire_con_in_stage5[74]), .outData_75(wire_con_in_stage5[75]), .outData_76(wire_con_in_stage5[76]), .outData_77(wire_con_in_stage5[77]), .outData_78(wire_con_in_stage5[78]), .outData_79(wire_con_in_stage5[79]), .outData_80(wire_con_in_stage5[80]), .outData_81(wire_con_in_stage5[81]), .outData_82(wire_con_in_stage5[82]), .outData_83(wire_con_in_stage5[83]), .outData_84(wire_con_in_stage5[84]), .outData_85(wire_con_in_stage5[85]), .outData_86(wire_con_in_stage5[86]), .outData_87(wire_con_in_stage5[87]), .outData_88(wire_con_in_stage5[88]), .outData_89(wire_con_in_stage5[89]), .outData_90(wire_con_in_stage5[90]), .outData_91(wire_con_in_stage5[91]), .outData_92(wire_con_in_stage5[92]), .outData_93(wire_con_in_stage5[93]), .outData_94(wire_con_in_stage5[94]), .outData_95(wire_con_in_stage5[95]), .outData_96(wire_con_in_stage5[96]), .outData_97(wire_con_in_stage5[97]), .outData_98(wire_con_in_stage5[98]), .outData_99(wire_con_in_stage5[99]), .outData_100(wire_con_in_stage5[100]), .outData_101(wire_con_in_stage5[101]), .outData_102(wire_con_in_stage5[102]), .outData_103(wire_con_in_stage5[103]), .outData_104(wire_con_in_stage5[104]), .outData_105(wire_con_in_stage5[105]), .outData_106(wire_con_in_stage5[106]), .outData_107(wire_con_in_stage5[107]), .outData_108(wire_con_in_stage5[108]), .outData_109(wire_con_in_stage5[109]), .outData_110(wire_con_in_stage5[110]), .outData_111(wire_con_in_stage5[111]), .outData_112(wire_con_in_stage5[112]), .outData_113(wire_con_in_stage5[113]), .outData_114(wire_con_in_stage5[114]), .outData_115(wire_con_in_stage5[115]), .outData_116(wire_con_in_stage5[116]), .outData_117(wire_con_in_stage5[117]), .outData_118(wire_con_in_stage5[118]), .outData_119(wire_con_in_stage5[119]), .outData_120(wire_con_in_stage5[120]), .outData_121(wire_con_in_stage5[121]), .outData_122(wire_con_in_stage5[122]), .outData_123(wire_con_in_stage5[123]), .outData_124(wire_con_in_stage5[124]), .outData_125(wire_con_in_stage5[125]), .outData_126(wire_con_in_stage5[126]), .outData_127(wire_con_in_stage5[127]), .outData_128(wire_con_in_stage5[128]), .outData_129(wire_con_in_stage5[129]), .outData_130(wire_con_in_stage5[130]), .outData_131(wire_con_in_stage5[131]), .outData_132(wire_con_in_stage5[132]), .outData_133(wire_con_in_stage5[133]), .outData_134(wire_con_in_stage5[134]), .outData_135(wire_con_in_stage5[135]), .outData_136(wire_con_in_stage5[136]), .outData_137(wire_con_in_stage5[137]), .outData_138(wire_con_in_stage5[138]), .outData_139(wire_con_in_stage5[139]), .outData_140(wire_con_in_stage5[140]), .outData_141(wire_con_in_stage5[141]), .outData_142(wire_con_in_stage5[142]), .outData_143(wire_con_in_stage5[143]), .outData_144(wire_con_in_stage5[144]), .outData_145(wire_con_in_stage5[145]), .outData_146(wire_con_in_stage5[146]), .outData_147(wire_con_in_stage5[147]), .outData_148(wire_con_in_stage5[148]), .outData_149(wire_con_in_stage5[149]), .outData_150(wire_con_in_stage5[150]), .outData_151(wire_con_in_stage5[151]), .outData_152(wire_con_in_stage5[152]), .outData_153(wire_con_in_stage5[153]), .outData_154(wire_con_in_stage5[154]), .outData_155(wire_con_in_stage5[155]), .outData_156(wire_con_in_stage5[156]), .outData_157(wire_con_in_stage5[157]), .outData_158(wire_con_in_stage5[158]), .outData_159(wire_con_in_stage5[159]), .outData_160(wire_con_in_stage5[160]), .outData_161(wire_con_in_stage5[161]), .outData_162(wire_con_in_stage5[162]), .outData_163(wire_con_in_stage5[163]), .outData_164(wire_con_in_stage5[164]), .outData_165(wire_con_in_stage5[165]), .outData_166(wire_con_in_stage5[166]), .outData_167(wire_con_in_stage5[167]), .outData_168(wire_con_in_stage5[168]), .outData_169(wire_con_in_stage5[169]), .outData_170(wire_con_in_stage5[170]), .outData_171(wire_con_in_stage5[171]), .outData_172(wire_con_in_stage5[172]), .outData_173(wire_con_in_stage5[173]), .outData_174(wire_con_in_stage5[174]), .outData_175(wire_con_in_stage5[175]), .outData_176(wire_con_in_stage5[176]), .outData_177(wire_con_in_stage5[177]), .outData_178(wire_con_in_stage5[178]), .outData_179(wire_con_in_stage5[179]), .outData_180(wire_con_in_stage5[180]), .outData_181(wire_con_in_stage5[181]), .outData_182(wire_con_in_stage5[182]), .outData_183(wire_con_in_stage5[183]), .outData_184(wire_con_in_stage5[184]), .outData_185(wire_con_in_stage5[185]), .outData_186(wire_con_in_stage5[186]), .outData_187(wire_con_in_stage5[187]), .outData_188(wire_con_in_stage5[188]), .outData_189(wire_con_in_stage5[189]), .outData_190(wire_con_in_stage5[190]), .outData_191(wire_con_in_stage5[191]), .outData_192(wire_con_in_stage5[192]), .outData_193(wire_con_in_stage5[193]), .outData_194(wire_con_in_stage5[194]), .outData_195(wire_con_in_stage5[195]), .outData_196(wire_con_in_stage5[196]), .outData_197(wire_con_in_stage5[197]), .outData_198(wire_con_in_stage5[198]), .outData_199(wire_con_in_stage5[199]), .outData_200(wire_con_in_stage5[200]), .outData_201(wire_con_in_stage5[201]), .outData_202(wire_con_in_stage5[202]), .outData_203(wire_con_in_stage5[203]), .outData_204(wire_con_in_stage5[204]), .outData_205(wire_con_in_stage5[205]), .outData_206(wire_con_in_stage5[206]), .outData_207(wire_con_in_stage5[207]), .outData_208(wire_con_in_stage5[208]), .outData_209(wire_con_in_stage5[209]), .outData_210(wire_con_in_stage5[210]), .outData_211(wire_con_in_stage5[211]), .outData_212(wire_con_in_stage5[212]), .outData_213(wire_con_in_stage5[213]), .outData_214(wire_con_in_stage5[214]), .outData_215(wire_con_in_stage5[215]), .outData_216(wire_con_in_stage5[216]), .outData_217(wire_con_in_stage5[217]), .outData_218(wire_con_in_stage5[218]), .outData_219(wire_con_in_stage5[219]), .outData_220(wire_con_in_stage5[220]), .outData_221(wire_con_in_stage5[221]), .outData_222(wire_con_in_stage5[222]), .outData_223(wire_con_in_stage5[223]), .outData_224(wire_con_in_stage5[224]), .outData_225(wire_con_in_stage5[225]), .outData_226(wire_con_in_stage5[226]), .outData_227(wire_con_in_stage5[227]), .outData_228(wire_con_in_stage5[228]), .outData_229(wire_con_in_stage5[229]), .outData_230(wire_con_in_stage5[230]), .outData_231(wire_con_in_stage5[231]), .outData_232(wire_con_in_stage5[232]), .outData_233(wire_con_in_stage5[233]), .outData_234(wire_con_in_stage5[234]), .outData_235(wire_con_in_stage5[235]), .outData_236(wire_con_in_stage5[236]), .outData_237(wire_con_in_stage5[237]), .outData_238(wire_con_in_stage5[238]), .outData_239(wire_con_in_stage5[239]), .outData_240(wire_con_in_stage5[240]), .outData_241(wire_con_in_stage5[241]), .outData_242(wire_con_in_stage5[242]), .outData_243(wire_con_in_stage5[243]), .outData_244(wire_con_in_stage5[244]), .outData_245(wire_con_in_stage5[245]), .outData_246(wire_con_in_stage5[246]), .outData_247(wire_con_in_stage5[247]), .outData_248(wire_con_in_stage5[248]), .outData_249(wire_con_in_stage5[249]), .outData_250(wire_con_in_stage5[250]), .outData_251(wire_con_in_stage5[251]), .outData_252(wire_con_in_stage5[252]), .outData_253(wire_con_in_stage5[253]), .outData_254(wire_con_in_stage5[254]), .outData_255(wire_con_in_stage5[255]), 
        .in_start(in_start_stage5), .out_start(con_in_start_stage5), .ctrl(wire_ctrl_stage5), .clk(clk), .rst(rst));
  
  wireCon_dp256_st5_L wire_stage_5(
        .inData_0(wire_con_in_stage5[0]), .inData_1(wire_con_in_stage5[1]), .inData_2(wire_con_in_stage5[2]), .inData_3(wire_con_in_stage5[3]), .inData_4(wire_con_in_stage5[4]), .inData_5(wire_con_in_stage5[5]), .inData_6(wire_con_in_stage5[6]), .inData_7(wire_con_in_stage5[7]), .inData_8(wire_con_in_stage5[8]), .inData_9(wire_con_in_stage5[9]), .inData_10(wire_con_in_stage5[10]), .inData_11(wire_con_in_stage5[11]), .inData_12(wire_con_in_stage5[12]), .inData_13(wire_con_in_stage5[13]), .inData_14(wire_con_in_stage5[14]), .inData_15(wire_con_in_stage5[15]), .inData_16(wire_con_in_stage5[16]), .inData_17(wire_con_in_stage5[17]), .inData_18(wire_con_in_stage5[18]), .inData_19(wire_con_in_stage5[19]), .inData_20(wire_con_in_stage5[20]), .inData_21(wire_con_in_stage5[21]), .inData_22(wire_con_in_stage5[22]), .inData_23(wire_con_in_stage5[23]), .inData_24(wire_con_in_stage5[24]), .inData_25(wire_con_in_stage5[25]), .inData_26(wire_con_in_stage5[26]), .inData_27(wire_con_in_stage5[27]), .inData_28(wire_con_in_stage5[28]), .inData_29(wire_con_in_stage5[29]), .inData_30(wire_con_in_stage5[30]), .inData_31(wire_con_in_stage5[31]), .inData_32(wire_con_in_stage5[32]), .inData_33(wire_con_in_stage5[33]), .inData_34(wire_con_in_stage5[34]), .inData_35(wire_con_in_stage5[35]), .inData_36(wire_con_in_stage5[36]), .inData_37(wire_con_in_stage5[37]), .inData_38(wire_con_in_stage5[38]), .inData_39(wire_con_in_stage5[39]), .inData_40(wire_con_in_stage5[40]), .inData_41(wire_con_in_stage5[41]), .inData_42(wire_con_in_stage5[42]), .inData_43(wire_con_in_stage5[43]), .inData_44(wire_con_in_stage5[44]), .inData_45(wire_con_in_stage5[45]), .inData_46(wire_con_in_stage5[46]), .inData_47(wire_con_in_stage5[47]), .inData_48(wire_con_in_stage5[48]), .inData_49(wire_con_in_stage5[49]), .inData_50(wire_con_in_stage5[50]), .inData_51(wire_con_in_stage5[51]), .inData_52(wire_con_in_stage5[52]), .inData_53(wire_con_in_stage5[53]), .inData_54(wire_con_in_stage5[54]), .inData_55(wire_con_in_stage5[55]), .inData_56(wire_con_in_stage5[56]), .inData_57(wire_con_in_stage5[57]), .inData_58(wire_con_in_stage5[58]), .inData_59(wire_con_in_stage5[59]), .inData_60(wire_con_in_stage5[60]), .inData_61(wire_con_in_stage5[61]), .inData_62(wire_con_in_stage5[62]), .inData_63(wire_con_in_stage5[63]), .inData_64(wire_con_in_stage5[64]), .inData_65(wire_con_in_stage5[65]), .inData_66(wire_con_in_stage5[66]), .inData_67(wire_con_in_stage5[67]), .inData_68(wire_con_in_stage5[68]), .inData_69(wire_con_in_stage5[69]), .inData_70(wire_con_in_stage5[70]), .inData_71(wire_con_in_stage5[71]), .inData_72(wire_con_in_stage5[72]), .inData_73(wire_con_in_stage5[73]), .inData_74(wire_con_in_stage5[74]), .inData_75(wire_con_in_stage5[75]), .inData_76(wire_con_in_stage5[76]), .inData_77(wire_con_in_stage5[77]), .inData_78(wire_con_in_stage5[78]), .inData_79(wire_con_in_stage5[79]), .inData_80(wire_con_in_stage5[80]), .inData_81(wire_con_in_stage5[81]), .inData_82(wire_con_in_stage5[82]), .inData_83(wire_con_in_stage5[83]), .inData_84(wire_con_in_stage5[84]), .inData_85(wire_con_in_stage5[85]), .inData_86(wire_con_in_stage5[86]), .inData_87(wire_con_in_stage5[87]), .inData_88(wire_con_in_stage5[88]), .inData_89(wire_con_in_stage5[89]), .inData_90(wire_con_in_stage5[90]), .inData_91(wire_con_in_stage5[91]), .inData_92(wire_con_in_stage5[92]), .inData_93(wire_con_in_stage5[93]), .inData_94(wire_con_in_stage5[94]), .inData_95(wire_con_in_stage5[95]), .inData_96(wire_con_in_stage5[96]), .inData_97(wire_con_in_stage5[97]), .inData_98(wire_con_in_stage5[98]), .inData_99(wire_con_in_stage5[99]), .inData_100(wire_con_in_stage5[100]), .inData_101(wire_con_in_stage5[101]), .inData_102(wire_con_in_stage5[102]), .inData_103(wire_con_in_stage5[103]), .inData_104(wire_con_in_stage5[104]), .inData_105(wire_con_in_stage5[105]), .inData_106(wire_con_in_stage5[106]), .inData_107(wire_con_in_stage5[107]), .inData_108(wire_con_in_stage5[108]), .inData_109(wire_con_in_stage5[109]), .inData_110(wire_con_in_stage5[110]), .inData_111(wire_con_in_stage5[111]), .inData_112(wire_con_in_stage5[112]), .inData_113(wire_con_in_stage5[113]), .inData_114(wire_con_in_stage5[114]), .inData_115(wire_con_in_stage5[115]), .inData_116(wire_con_in_stage5[116]), .inData_117(wire_con_in_stage5[117]), .inData_118(wire_con_in_stage5[118]), .inData_119(wire_con_in_stage5[119]), .inData_120(wire_con_in_stage5[120]), .inData_121(wire_con_in_stage5[121]), .inData_122(wire_con_in_stage5[122]), .inData_123(wire_con_in_stage5[123]), .inData_124(wire_con_in_stage5[124]), .inData_125(wire_con_in_stage5[125]), .inData_126(wire_con_in_stage5[126]), .inData_127(wire_con_in_stage5[127]), .inData_128(wire_con_in_stage5[128]), .inData_129(wire_con_in_stage5[129]), .inData_130(wire_con_in_stage5[130]), .inData_131(wire_con_in_stage5[131]), .inData_132(wire_con_in_stage5[132]), .inData_133(wire_con_in_stage5[133]), .inData_134(wire_con_in_stage5[134]), .inData_135(wire_con_in_stage5[135]), .inData_136(wire_con_in_stage5[136]), .inData_137(wire_con_in_stage5[137]), .inData_138(wire_con_in_stage5[138]), .inData_139(wire_con_in_stage5[139]), .inData_140(wire_con_in_stage5[140]), .inData_141(wire_con_in_stage5[141]), .inData_142(wire_con_in_stage5[142]), .inData_143(wire_con_in_stage5[143]), .inData_144(wire_con_in_stage5[144]), .inData_145(wire_con_in_stage5[145]), .inData_146(wire_con_in_stage5[146]), .inData_147(wire_con_in_stage5[147]), .inData_148(wire_con_in_stage5[148]), .inData_149(wire_con_in_stage5[149]), .inData_150(wire_con_in_stage5[150]), .inData_151(wire_con_in_stage5[151]), .inData_152(wire_con_in_stage5[152]), .inData_153(wire_con_in_stage5[153]), .inData_154(wire_con_in_stage5[154]), .inData_155(wire_con_in_stage5[155]), .inData_156(wire_con_in_stage5[156]), .inData_157(wire_con_in_stage5[157]), .inData_158(wire_con_in_stage5[158]), .inData_159(wire_con_in_stage5[159]), .inData_160(wire_con_in_stage5[160]), .inData_161(wire_con_in_stage5[161]), .inData_162(wire_con_in_stage5[162]), .inData_163(wire_con_in_stage5[163]), .inData_164(wire_con_in_stage5[164]), .inData_165(wire_con_in_stage5[165]), .inData_166(wire_con_in_stage5[166]), .inData_167(wire_con_in_stage5[167]), .inData_168(wire_con_in_stage5[168]), .inData_169(wire_con_in_stage5[169]), .inData_170(wire_con_in_stage5[170]), .inData_171(wire_con_in_stage5[171]), .inData_172(wire_con_in_stage5[172]), .inData_173(wire_con_in_stage5[173]), .inData_174(wire_con_in_stage5[174]), .inData_175(wire_con_in_stage5[175]), .inData_176(wire_con_in_stage5[176]), .inData_177(wire_con_in_stage5[177]), .inData_178(wire_con_in_stage5[178]), .inData_179(wire_con_in_stage5[179]), .inData_180(wire_con_in_stage5[180]), .inData_181(wire_con_in_stage5[181]), .inData_182(wire_con_in_stage5[182]), .inData_183(wire_con_in_stage5[183]), .inData_184(wire_con_in_stage5[184]), .inData_185(wire_con_in_stage5[185]), .inData_186(wire_con_in_stage5[186]), .inData_187(wire_con_in_stage5[187]), .inData_188(wire_con_in_stage5[188]), .inData_189(wire_con_in_stage5[189]), .inData_190(wire_con_in_stage5[190]), .inData_191(wire_con_in_stage5[191]), .inData_192(wire_con_in_stage5[192]), .inData_193(wire_con_in_stage5[193]), .inData_194(wire_con_in_stage5[194]), .inData_195(wire_con_in_stage5[195]), .inData_196(wire_con_in_stage5[196]), .inData_197(wire_con_in_stage5[197]), .inData_198(wire_con_in_stage5[198]), .inData_199(wire_con_in_stage5[199]), .inData_200(wire_con_in_stage5[200]), .inData_201(wire_con_in_stage5[201]), .inData_202(wire_con_in_stage5[202]), .inData_203(wire_con_in_stage5[203]), .inData_204(wire_con_in_stage5[204]), .inData_205(wire_con_in_stage5[205]), .inData_206(wire_con_in_stage5[206]), .inData_207(wire_con_in_stage5[207]), .inData_208(wire_con_in_stage5[208]), .inData_209(wire_con_in_stage5[209]), .inData_210(wire_con_in_stage5[210]), .inData_211(wire_con_in_stage5[211]), .inData_212(wire_con_in_stage5[212]), .inData_213(wire_con_in_stage5[213]), .inData_214(wire_con_in_stage5[214]), .inData_215(wire_con_in_stage5[215]), .inData_216(wire_con_in_stage5[216]), .inData_217(wire_con_in_stage5[217]), .inData_218(wire_con_in_stage5[218]), .inData_219(wire_con_in_stage5[219]), .inData_220(wire_con_in_stage5[220]), .inData_221(wire_con_in_stage5[221]), .inData_222(wire_con_in_stage5[222]), .inData_223(wire_con_in_stage5[223]), .inData_224(wire_con_in_stage5[224]), .inData_225(wire_con_in_stage5[225]), .inData_226(wire_con_in_stage5[226]), .inData_227(wire_con_in_stage5[227]), .inData_228(wire_con_in_stage5[228]), .inData_229(wire_con_in_stage5[229]), .inData_230(wire_con_in_stage5[230]), .inData_231(wire_con_in_stage5[231]), .inData_232(wire_con_in_stage5[232]), .inData_233(wire_con_in_stage5[233]), .inData_234(wire_con_in_stage5[234]), .inData_235(wire_con_in_stage5[235]), .inData_236(wire_con_in_stage5[236]), .inData_237(wire_con_in_stage5[237]), .inData_238(wire_con_in_stage5[238]), .inData_239(wire_con_in_stage5[239]), .inData_240(wire_con_in_stage5[240]), .inData_241(wire_con_in_stage5[241]), .inData_242(wire_con_in_stage5[242]), .inData_243(wire_con_in_stage5[243]), .inData_244(wire_con_in_stage5[244]), .inData_245(wire_con_in_stage5[245]), .inData_246(wire_con_in_stage5[246]), .inData_247(wire_con_in_stage5[247]), .inData_248(wire_con_in_stage5[248]), .inData_249(wire_con_in_stage5[249]), .inData_250(wire_con_in_stage5[250]), .inData_251(wire_con_in_stage5[251]), .inData_252(wire_con_in_stage5[252]), .inData_253(wire_con_in_stage5[253]), .inData_254(wire_con_in_stage5[254]), .inData_255(wire_con_in_stage5[255]), 
        .outData_0(wire_con_out_stage5[0]), .outData_1(wire_con_out_stage5[1]), .outData_2(wire_con_out_stage5[2]), .outData_3(wire_con_out_stage5[3]), .outData_4(wire_con_out_stage5[4]), .outData_5(wire_con_out_stage5[5]), .outData_6(wire_con_out_stage5[6]), .outData_7(wire_con_out_stage5[7]), .outData_8(wire_con_out_stage5[8]), .outData_9(wire_con_out_stage5[9]), .outData_10(wire_con_out_stage5[10]), .outData_11(wire_con_out_stage5[11]), .outData_12(wire_con_out_stage5[12]), .outData_13(wire_con_out_stage5[13]), .outData_14(wire_con_out_stage5[14]), .outData_15(wire_con_out_stage5[15]), .outData_16(wire_con_out_stage5[16]), .outData_17(wire_con_out_stage5[17]), .outData_18(wire_con_out_stage5[18]), .outData_19(wire_con_out_stage5[19]), .outData_20(wire_con_out_stage5[20]), .outData_21(wire_con_out_stage5[21]), .outData_22(wire_con_out_stage5[22]), .outData_23(wire_con_out_stage5[23]), .outData_24(wire_con_out_stage5[24]), .outData_25(wire_con_out_stage5[25]), .outData_26(wire_con_out_stage5[26]), .outData_27(wire_con_out_stage5[27]), .outData_28(wire_con_out_stage5[28]), .outData_29(wire_con_out_stage5[29]), .outData_30(wire_con_out_stage5[30]), .outData_31(wire_con_out_stage5[31]), .outData_32(wire_con_out_stage5[32]), .outData_33(wire_con_out_stage5[33]), .outData_34(wire_con_out_stage5[34]), .outData_35(wire_con_out_stage5[35]), .outData_36(wire_con_out_stage5[36]), .outData_37(wire_con_out_stage5[37]), .outData_38(wire_con_out_stage5[38]), .outData_39(wire_con_out_stage5[39]), .outData_40(wire_con_out_stage5[40]), .outData_41(wire_con_out_stage5[41]), .outData_42(wire_con_out_stage5[42]), .outData_43(wire_con_out_stage5[43]), .outData_44(wire_con_out_stage5[44]), .outData_45(wire_con_out_stage5[45]), .outData_46(wire_con_out_stage5[46]), .outData_47(wire_con_out_stage5[47]), .outData_48(wire_con_out_stage5[48]), .outData_49(wire_con_out_stage5[49]), .outData_50(wire_con_out_stage5[50]), .outData_51(wire_con_out_stage5[51]), .outData_52(wire_con_out_stage5[52]), .outData_53(wire_con_out_stage5[53]), .outData_54(wire_con_out_stage5[54]), .outData_55(wire_con_out_stage5[55]), .outData_56(wire_con_out_stage5[56]), .outData_57(wire_con_out_stage5[57]), .outData_58(wire_con_out_stage5[58]), .outData_59(wire_con_out_stage5[59]), .outData_60(wire_con_out_stage5[60]), .outData_61(wire_con_out_stage5[61]), .outData_62(wire_con_out_stage5[62]), .outData_63(wire_con_out_stage5[63]), .outData_64(wire_con_out_stage5[64]), .outData_65(wire_con_out_stage5[65]), .outData_66(wire_con_out_stage5[66]), .outData_67(wire_con_out_stage5[67]), .outData_68(wire_con_out_stage5[68]), .outData_69(wire_con_out_stage5[69]), .outData_70(wire_con_out_stage5[70]), .outData_71(wire_con_out_stage5[71]), .outData_72(wire_con_out_stage5[72]), .outData_73(wire_con_out_stage5[73]), .outData_74(wire_con_out_stage5[74]), .outData_75(wire_con_out_stage5[75]), .outData_76(wire_con_out_stage5[76]), .outData_77(wire_con_out_stage5[77]), .outData_78(wire_con_out_stage5[78]), .outData_79(wire_con_out_stage5[79]), .outData_80(wire_con_out_stage5[80]), .outData_81(wire_con_out_stage5[81]), .outData_82(wire_con_out_stage5[82]), .outData_83(wire_con_out_stage5[83]), .outData_84(wire_con_out_stage5[84]), .outData_85(wire_con_out_stage5[85]), .outData_86(wire_con_out_stage5[86]), .outData_87(wire_con_out_stage5[87]), .outData_88(wire_con_out_stage5[88]), .outData_89(wire_con_out_stage5[89]), .outData_90(wire_con_out_stage5[90]), .outData_91(wire_con_out_stage5[91]), .outData_92(wire_con_out_stage5[92]), .outData_93(wire_con_out_stage5[93]), .outData_94(wire_con_out_stage5[94]), .outData_95(wire_con_out_stage5[95]), .outData_96(wire_con_out_stage5[96]), .outData_97(wire_con_out_stage5[97]), .outData_98(wire_con_out_stage5[98]), .outData_99(wire_con_out_stage5[99]), .outData_100(wire_con_out_stage5[100]), .outData_101(wire_con_out_stage5[101]), .outData_102(wire_con_out_stage5[102]), .outData_103(wire_con_out_stage5[103]), .outData_104(wire_con_out_stage5[104]), .outData_105(wire_con_out_stage5[105]), .outData_106(wire_con_out_stage5[106]), .outData_107(wire_con_out_stage5[107]), .outData_108(wire_con_out_stage5[108]), .outData_109(wire_con_out_stage5[109]), .outData_110(wire_con_out_stage5[110]), .outData_111(wire_con_out_stage5[111]), .outData_112(wire_con_out_stage5[112]), .outData_113(wire_con_out_stage5[113]), .outData_114(wire_con_out_stage5[114]), .outData_115(wire_con_out_stage5[115]), .outData_116(wire_con_out_stage5[116]), .outData_117(wire_con_out_stage5[117]), .outData_118(wire_con_out_stage5[118]), .outData_119(wire_con_out_stage5[119]), .outData_120(wire_con_out_stage5[120]), .outData_121(wire_con_out_stage5[121]), .outData_122(wire_con_out_stage5[122]), .outData_123(wire_con_out_stage5[123]), .outData_124(wire_con_out_stage5[124]), .outData_125(wire_con_out_stage5[125]), .outData_126(wire_con_out_stage5[126]), .outData_127(wire_con_out_stage5[127]), .outData_128(wire_con_out_stage5[128]), .outData_129(wire_con_out_stage5[129]), .outData_130(wire_con_out_stage5[130]), .outData_131(wire_con_out_stage5[131]), .outData_132(wire_con_out_stage5[132]), .outData_133(wire_con_out_stage5[133]), .outData_134(wire_con_out_stage5[134]), .outData_135(wire_con_out_stage5[135]), .outData_136(wire_con_out_stage5[136]), .outData_137(wire_con_out_stage5[137]), .outData_138(wire_con_out_stage5[138]), .outData_139(wire_con_out_stage5[139]), .outData_140(wire_con_out_stage5[140]), .outData_141(wire_con_out_stage5[141]), .outData_142(wire_con_out_stage5[142]), .outData_143(wire_con_out_stage5[143]), .outData_144(wire_con_out_stage5[144]), .outData_145(wire_con_out_stage5[145]), .outData_146(wire_con_out_stage5[146]), .outData_147(wire_con_out_stage5[147]), .outData_148(wire_con_out_stage5[148]), .outData_149(wire_con_out_stage5[149]), .outData_150(wire_con_out_stage5[150]), .outData_151(wire_con_out_stage5[151]), .outData_152(wire_con_out_stage5[152]), .outData_153(wire_con_out_stage5[153]), .outData_154(wire_con_out_stage5[154]), .outData_155(wire_con_out_stage5[155]), .outData_156(wire_con_out_stage5[156]), .outData_157(wire_con_out_stage5[157]), .outData_158(wire_con_out_stage5[158]), .outData_159(wire_con_out_stage5[159]), .outData_160(wire_con_out_stage5[160]), .outData_161(wire_con_out_stage5[161]), .outData_162(wire_con_out_stage5[162]), .outData_163(wire_con_out_stage5[163]), .outData_164(wire_con_out_stage5[164]), .outData_165(wire_con_out_stage5[165]), .outData_166(wire_con_out_stage5[166]), .outData_167(wire_con_out_stage5[167]), .outData_168(wire_con_out_stage5[168]), .outData_169(wire_con_out_stage5[169]), .outData_170(wire_con_out_stage5[170]), .outData_171(wire_con_out_stage5[171]), .outData_172(wire_con_out_stage5[172]), .outData_173(wire_con_out_stage5[173]), .outData_174(wire_con_out_stage5[174]), .outData_175(wire_con_out_stage5[175]), .outData_176(wire_con_out_stage5[176]), .outData_177(wire_con_out_stage5[177]), .outData_178(wire_con_out_stage5[178]), .outData_179(wire_con_out_stage5[179]), .outData_180(wire_con_out_stage5[180]), .outData_181(wire_con_out_stage5[181]), .outData_182(wire_con_out_stage5[182]), .outData_183(wire_con_out_stage5[183]), .outData_184(wire_con_out_stage5[184]), .outData_185(wire_con_out_stage5[185]), .outData_186(wire_con_out_stage5[186]), .outData_187(wire_con_out_stage5[187]), .outData_188(wire_con_out_stage5[188]), .outData_189(wire_con_out_stage5[189]), .outData_190(wire_con_out_stage5[190]), .outData_191(wire_con_out_stage5[191]), .outData_192(wire_con_out_stage5[192]), .outData_193(wire_con_out_stage5[193]), .outData_194(wire_con_out_stage5[194]), .outData_195(wire_con_out_stage5[195]), .outData_196(wire_con_out_stage5[196]), .outData_197(wire_con_out_stage5[197]), .outData_198(wire_con_out_stage5[198]), .outData_199(wire_con_out_stage5[199]), .outData_200(wire_con_out_stage5[200]), .outData_201(wire_con_out_stage5[201]), .outData_202(wire_con_out_stage5[202]), .outData_203(wire_con_out_stage5[203]), .outData_204(wire_con_out_stage5[204]), .outData_205(wire_con_out_stage5[205]), .outData_206(wire_con_out_stage5[206]), .outData_207(wire_con_out_stage5[207]), .outData_208(wire_con_out_stage5[208]), .outData_209(wire_con_out_stage5[209]), .outData_210(wire_con_out_stage5[210]), .outData_211(wire_con_out_stage5[211]), .outData_212(wire_con_out_stage5[212]), .outData_213(wire_con_out_stage5[213]), .outData_214(wire_con_out_stage5[214]), .outData_215(wire_con_out_stage5[215]), .outData_216(wire_con_out_stage5[216]), .outData_217(wire_con_out_stage5[217]), .outData_218(wire_con_out_stage5[218]), .outData_219(wire_con_out_stage5[219]), .outData_220(wire_con_out_stage5[220]), .outData_221(wire_con_out_stage5[221]), .outData_222(wire_con_out_stage5[222]), .outData_223(wire_con_out_stage5[223]), .outData_224(wire_con_out_stage5[224]), .outData_225(wire_con_out_stage5[225]), .outData_226(wire_con_out_stage5[226]), .outData_227(wire_con_out_stage5[227]), .outData_228(wire_con_out_stage5[228]), .outData_229(wire_con_out_stage5[229]), .outData_230(wire_con_out_stage5[230]), .outData_231(wire_con_out_stage5[231]), .outData_232(wire_con_out_stage5[232]), .outData_233(wire_con_out_stage5[233]), .outData_234(wire_con_out_stage5[234]), .outData_235(wire_con_out_stage5[235]), .outData_236(wire_con_out_stage5[236]), .outData_237(wire_con_out_stage5[237]), .outData_238(wire_con_out_stage5[238]), .outData_239(wire_con_out_stage5[239]), .outData_240(wire_con_out_stage5[240]), .outData_241(wire_con_out_stage5[241]), .outData_242(wire_con_out_stage5[242]), .outData_243(wire_con_out_stage5[243]), .outData_244(wire_con_out_stage5[244]), .outData_245(wire_con_out_stage5[245]), .outData_246(wire_con_out_stage5[246]), .outData_247(wire_con_out_stage5[247]), .outData_248(wire_con_out_stage5[248]), .outData_249(wire_con_out_stage5[249]), .outData_250(wire_con_out_stage5[250]), .outData_251(wire_con_out_stage5[251]), .outData_252(wire_con_out_stage5[252]), .outData_253(wire_con_out_stage5[253]), .outData_254(wire_con_out_stage5[254]), .outData_255(wire_con_out_stage5[255]), 
        .in_start(con_in_start_stage5), .out_start(in_start_stage6), .clk(clk), .rst(rst)); 

  
  assign wire_ctrl_stage5[0] = counter_w[2]; 
  assign wire_ctrl_stage5[1] = counter_w[2]; 
  assign wire_ctrl_stage5[2] = counter_w[2]; 
  assign wire_ctrl_stage5[3] = counter_w[2]; 
  assign wire_ctrl_stage5[4] = counter_w[2]; 
  assign wire_ctrl_stage5[5] = counter_w[2]; 
  assign wire_ctrl_stage5[6] = counter_w[2]; 
  assign wire_ctrl_stage5[7] = counter_w[2]; 
  assign wire_ctrl_stage5[8] = counter_w[2]; 
  assign wire_ctrl_stage5[9] = counter_w[2]; 
  assign wire_ctrl_stage5[10] = counter_w[2]; 
  assign wire_ctrl_stage5[11] = counter_w[2]; 
  assign wire_ctrl_stage5[12] = counter_w[2]; 
  assign wire_ctrl_stage5[13] = counter_w[2]; 
  assign wire_ctrl_stage5[14] = counter_w[2]; 
  assign wire_ctrl_stage5[15] = counter_w[2]; 
  assign wire_ctrl_stage5[16] = counter_w[2]; 
  assign wire_ctrl_stage5[17] = counter_w[2]; 
  assign wire_ctrl_stage5[18] = counter_w[2]; 
  assign wire_ctrl_stage5[19] = counter_w[2]; 
  assign wire_ctrl_stage5[20] = counter_w[2]; 
  assign wire_ctrl_stage5[21] = counter_w[2]; 
  assign wire_ctrl_stage5[22] = counter_w[2]; 
  assign wire_ctrl_stage5[23] = counter_w[2]; 
  assign wire_ctrl_stage5[24] = counter_w[2]; 
  assign wire_ctrl_stage5[25] = counter_w[2]; 
  assign wire_ctrl_stage5[26] = counter_w[2]; 
  assign wire_ctrl_stage5[27] = counter_w[2]; 
  assign wire_ctrl_stage5[28] = counter_w[2]; 
  assign wire_ctrl_stage5[29] = counter_w[2]; 
  assign wire_ctrl_stage5[30] = counter_w[2]; 
  assign wire_ctrl_stage5[31] = counter_w[2]; 
  assign wire_ctrl_stage5[32] = counter_w[2]; 
  assign wire_ctrl_stage5[33] = counter_w[2]; 
  assign wire_ctrl_stage5[34] = counter_w[2]; 
  assign wire_ctrl_stage5[35] = counter_w[2]; 
  assign wire_ctrl_stage5[36] = counter_w[2]; 
  assign wire_ctrl_stage5[37] = counter_w[2]; 
  assign wire_ctrl_stage5[38] = counter_w[2]; 
  assign wire_ctrl_stage5[39] = counter_w[2]; 
  assign wire_ctrl_stage5[40] = counter_w[2]; 
  assign wire_ctrl_stage5[41] = counter_w[2]; 
  assign wire_ctrl_stage5[42] = counter_w[2]; 
  assign wire_ctrl_stage5[43] = counter_w[2]; 
  assign wire_ctrl_stage5[44] = counter_w[2]; 
  assign wire_ctrl_stage5[45] = counter_w[2]; 
  assign wire_ctrl_stage5[46] = counter_w[2]; 
  assign wire_ctrl_stage5[47] = counter_w[2]; 
  assign wire_ctrl_stage5[48] = counter_w[2]; 
  assign wire_ctrl_stage5[49] = counter_w[2]; 
  assign wire_ctrl_stage5[50] = counter_w[2]; 
  assign wire_ctrl_stage5[51] = counter_w[2]; 
  assign wire_ctrl_stage5[52] = counter_w[2]; 
  assign wire_ctrl_stage5[53] = counter_w[2]; 
  assign wire_ctrl_stage5[54] = counter_w[2]; 
  assign wire_ctrl_stage5[55] = counter_w[2]; 
  assign wire_ctrl_stage5[56] = counter_w[2]; 
  assign wire_ctrl_stage5[57] = counter_w[2]; 
  assign wire_ctrl_stage5[58] = counter_w[2]; 
  assign wire_ctrl_stage5[59] = counter_w[2]; 
  assign wire_ctrl_stage5[60] = counter_w[2]; 
  assign wire_ctrl_stage5[61] = counter_w[2]; 
  assign wire_ctrl_stage5[62] = counter_w[2]; 
  assign wire_ctrl_stage5[63] = counter_w[2]; 
  assign wire_ctrl_stage5[64] = counter_w[2]; 
  assign wire_ctrl_stage5[65] = counter_w[2]; 
  assign wire_ctrl_stage5[66] = counter_w[2]; 
  assign wire_ctrl_stage5[67] = counter_w[2]; 
  assign wire_ctrl_stage5[68] = counter_w[2]; 
  assign wire_ctrl_stage5[69] = counter_w[2]; 
  assign wire_ctrl_stage5[70] = counter_w[2]; 
  assign wire_ctrl_stage5[71] = counter_w[2]; 
  assign wire_ctrl_stage5[72] = counter_w[2]; 
  assign wire_ctrl_stage5[73] = counter_w[2]; 
  assign wire_ctrl_stage5[74] = counter_w[2]; 
  assign wire_ctrl_stage5[75] = counter_w[2]; 
  assign wire_ctrl_stage5[76] = counter_w[2]; 
  assign wire_ctrl_stage5[77] = counter_w[2]; 
  assign wire_ctrl_stage5[78] = counter_w[2]; 
  assign wire_ctrl_stage5[79] = counter_w[2]; 
  assign wire_ctrl_stage5[80] = counter_w[2]; 
  assign wire_ctrl_stage5[81] = counter_w[2]; 
  assign wire_ctrl_stage5[82] = counter_w[2]; 
  assign wire_ctrl_stage5[83] = counter_w[2]; 
  assign wire_ctrl_stage5[84] = counter_w[2]; 
  assign wire_ctrl_stage5[85] = counter_w[2]; 
  assign wire_ctrl_stage5[86] = counter_w[2]; 
  assign wire_ctrl_stage5[87] = counter_w[2]; 
  assign wire_ctrl_stage5[88] = counter_w[2]; 
  assign wire_ctrl_stage5[89] = counter_w[2]; 
  assign wire_ctrl_stage5[90] = counter_w[2]; 
  assign wire_ctrl_stage5[91] = counter_w[2]; 
  assign wire_ctrl_stage5[92] = counter_w[2]; 
  assign wire_ctrl_stage5[93] = counter_w[2]; 
  assign wire_ctrl_stage5[94] = counter_w[2]; 
  assign wire_ctrl_stage5[95] = counter_w[2]; 
  assign wire_ctrl_stage5[96] = counter_w[2]; 
  assign wire_ctrl_stage5[97] = counter_w[2]; 
  assign wire_ctrl_stage5[98] = counter_w[2]; 
  assign wire_ctrl_stage5[99] = counter_w[2]; 
  assign wire_ctrl_stage5[100] = counter_w[2]; 
  assign wire_ctrl_stage5[101] = counter_w[2]; 
  assign wire_ctrl_stage5[102] = counter_w[2]; 
  assign wire_ctrl_stage5[103] = counter_w[2]; 
  assign wire_ctrl_stage5[104] = counter_w[2]; 
  assign wire_ctrl_stage5[105] = counter_w[2]; 
  assign wire_ctrl_stage5[106] = counter_w[2]; 
  assign wire_ctrl_stage5[107] = counter_w[2]; 
  assign wire_ctrl_stage5[108] = counter_w[2]; 
  assign wire_ctrl_stage5[109] = counter_w[2]; 
  assign wire_ctrl_stage5[110] = counter_w[2]; 
  assign wire_ctrl_stage5[111] = counter_w[2]; 
  assign wire_ctrl_stage5[112] = counter_w[2]; 
  assign wire_ctrl_stage5[113] = counter_w[2]; 
  assign wire_ctrl_stage5[114] = counter_w[2]; 
  assign wire_ctrl_stage5[115] = counter_w[2]; 
  assign wire_ctrl_stage5[116] = counter_w[2]; 
  assign wire_ctrl_stage5[117] = counter_w[2]; 
  assign wire_ctrl_stage5[118] = counter_w[2]; 
  assign wire_ctrl_stage5[119] = counter_w[2]; 
  assign wire_ctrl_stage5[120] = counter_w[2]; 
  assign wire_ctrl_stage5[121] = counter_w[2]; 
  assign wire_ctrl_stage5[122] = counter_w[2]; 
  assign wire_ctrl_stage5[123] = counter_w[2]; 
  assign wire_ctrl_stage5[124] = counter_w[2]; 
  assign wire_ctrl_stage5[125] = counter_w[2]; 
  assign wire_ctrl_stage5[126] = counter_w[2]; 
  assign wire_ctrl_stage5[127] = counter_w[2]; 
  wire [DATA_WIDTH-1:0] wire_con_in_stage6[255:0];
  wire [DATA_WIDTH-1:0] wire_con_out_stage6[255:0];
  wire [127:0] wire_ctrl_stage6;

  switches_stage_st6_0_L switch_stage_6(
        .inData_0(wire_con_out_stage5[0]), .inData_1(wire_con_out_stage5[1]), .inData_2(wire_con_out_stage5[2]), .inData_3(wire_con_out_stage5[3]), .inData_4(wire_con_out_stage5[4]), .inData_5(wire_con_out_stage5[5]), .inData_6(wire_con_out_stage5[6]), .inData_7(wire_con_out_stage5[7]), .inData_8(wire_con_out_stage5[8]), .inData_9(wire_con_out_stage5[9]), .inData_10(wire_con_out_stage5[10]), .inData_11(wire_con_out_stage5[11]), .inData_12(wire_con_out_stage5[12]), .inData_13(wire_con_out_stage5[13]), .inData_14(wire_con_out_stage5[14]), .inData_15(wire_con_out_stage5[15]), .inData_16(wire_con_out_stage5[16]), .inData_17(wire_con_out_stage5[17]), .inData_18(wire_con_out_stage5[18]), .inData_19(wire_con_out_stage5[19]), .inData_20(wire_con_out_stage5[20]), .inData_21(wire_con_out_stage5[21]), .inData_22(wire_con_out_stage5[22]), .inData_23(wire_con_out_stage5[23]), .inData_24(wire_con_out_stage5[24]), .inData_25(wire_con_out_stage5[25]), .inData_26(wire_con_out_stage5[26]), .inData_27(wire_con_out_stage5[27]), .inData_28(wire_con_out_stage5[28]), .inData_29(wire_con_out_stage5[29]), .inData_30(wire_con_out_stage5[30]), .inData_31(wire_con_out_stage5[31]), .inData_32(wire_con_out_stage5[32]), .inData_33(wire_con_out_stage5[33]), .inData_34(wire_con_out_stage5[34]), .inData_35(wire_con_out_stage5[35]), .inData_36(wire_con_out_stage5[36]), .inData_37(wire_con_out_stage5[37]), .inData_38(wire_con_out_stage5[38]), .inData_39(wire_con_out_stage5[39]), .inData_40(wire_con_out_stage5[40]), .inData_41(wire_con_out_stage5[41]), .inData_42(wire_con_out_stage5[42]), .inData_43(wire_con_out_stage5[43]), .inData_44(wire_con_out_stage5[44]), .inData_45(wire_con_out_stage5[45]), .inData_46(wire_con_out_stage5[46]), .inData_47(wire_con_out_stage5[47]), .inData_48(wire_con_out_stage5[48]), .inData_49(wire_con_out_stage5[49]), .inData_50(wire_con_out_stage5[50]), .inData_51(wire_con_out_stage5[51]), .inData_52(wire_con_out_stage5[52]), .inData_53(wire_con_out_stage5[53]), .inData_54(wire_con_out_stage5[54]), .inData_55(wire_con_out_stage5[55]), .inData_56(wire_con_out_stage5[56]), .inData_57(wire_con_out_stage5[57]), .inData_58(wire_con_out_stage5[58]), .inData_59(wire_con_out_stage5[59]), .inData_60(wire_con_out_stage5[60]), .inData_61(wire_con_out_stage5[61]), .inData_62(wire_con_out_stage5[62]), .inData_63(wire_con_out_stage5[63]), .inData_64(wire_con_out_stage5[64]), .inData_65(wire_con_out_stage5[65]), .inData_66(wire_con_out_stage5[66]), .inData_67(wire_con_out_stage5[67]), .inData_68(wire_con_out_stage5[68]), .inData_69(wire_con_out_stage5[69]), .inData_70(wire_con_out_stage5[70]), .inData_71(wire_con_out_stage5[71]), .inData_72(wire_con_out_stage5[72]), .inData_73(wire_con_out_stage5[73]), .inData_74(wire_con_out_stage5[74]), .inData_75(wire_con_out_stage5[75]), .inData_76(wire_con_out_stage5[76]), .inData_77(wire_con_out_stage5[77]), .inData_78(wire_con_out_stage5[78]), .inData_79(wire_con_out_stage5[79]), .inData_80(wire_con_out_stage5[80]), .inData_81(wire_con_out_stage5[81]), .inData_82(wire_con_out_stage5[82]), .inData_83(wire_con_out_stage5[83]), .inData_84(wire_con_out_stage5[84]), .inData_85(wire_con_out_stage5[85]), .inData_86(wire_con_out_stage5[86]), .inData_87(wire_con_out_stage5[87]), .inData_88(wire_con_out_stage5[88]), .inData_89(wire_con_out_stage5[89]), .inData_90(wire_con_out_stage5[90]), .inData_91(wire_con_out_stage5[91]), .inData_92(wire_con_out_stage5[92]), .inData_93(wire_con_out_stage5[93]), .inData_94(wire_con_out_stage5[94]), .inData_95(wire_con_out_stage5[95]), .inData_96(wire_con_out_stage5[96]), .inData_97(wire_con_out_stage5[97]), .inData_98(wire_con_out_stage5[98]), .inData_99(wire_con_out_stage5[99]), .inData_100(wire_con_out_stage5[100]), .inData_101(wire_con_out_stage5[101]), .inData_102(wire_con_out_stage5[102]), .inData_103(wire_con_out_stage5[103]), .inData_104(wire_con_out_stage5[104]), .inData_105(wire_con_out_stage5[105]), .inData_106(wire_con_out_stage5[106]), .inData_107(wire_con_out_stage5[107]), .inData_108(wire_con_out_stage5[108]), .inData_109(wire_con_out_stage5[109]), .inData_110(wire_con_out_stage5[110]), .inData_111(wire_con_out_stage5[111]), .inData_112(wire_con_out_stage5[112]), .inData_113(wire_con_out_stage5[113]), .inData_114(wire_con_out_stage5[114]), .inData_115(wire_con_out_stage5[115]), .inData_116(wire_con_out_stage5[116]), .inData_117(wire_con_out_stage5[117]), .inData_118(wire_con_out_stage5[118]), .inData_119(wire_con_out_stage5[119]), .inData_120(wire_con_out_stage5[120]), .inData_121(wire_con_out_stage5[121]), .inData_122(wire_con_out_stage5[122]), .inData_123(wire_con_out_stage5[123]), .inData_124(wire_con_out_stage5[124]), .inData_125(wire_con_out_stage5[125]), .inData_126(wire_con_out_stage5[126]), .inData_127(wire_con_out_stage5[127]), .inData_128(wire_con_out_stage5[128]), .inData_129(wire_con_out_stage5[129]), .inData_130(wire_con_out_stage5[130]), .inData_131(wire_con_out_stage5[131]), .inData_132(wire_con_out_stage5[132]), .inData_133(wire_con_out_stage5[133]), .inData_134(wire_con_out_stage5[134]), .inData_135(wire_con_out_stage5[135]), .inData_136(wire_con_out_stage5[136]), .inData_137(wire_con_out_stage5[137]), .inData_138(wire_con_out_stage5[138]), .inData_139(wire_con_out_stage5[139]), .inData_140(wire_con_out_stage5[140]), .inData_141(wire_con_out_stage5[141]), .inData_142(wire_con_out_stage5[142]), .inData_143(wire_con_out_stage5[143]), .inData_144(wire_con_out_stage5[144]), .inData_145(wire_con_out_stage5[145]), .inData_146(wire_con_out_stage5[146]), .inData_147(wire_con_out_stage5[147]), .inData_148(wire_con_out_stage5[148]), .inData_149(wire_con_out_stage5[149]), .inData_150(wire_con_out_stage5[150]), .inData_151(wire_con_out_stage5[151]), .inData_152(wire_con_out_stage5[152]), .inData_153(wire_con_out_stage5[153]), .inData_154(wire_con_out_stage5[154]), .inData_155(wire_con_out_stage5[155]), .inData_156(wire_con_out_stage5[156]), .inData_157(wire_con_out_stage5[157]), .inData_158(wire_con_out_stage5[158]), .inData_159(wire_con_out_stage5[159]), .inData_160(wire_con_out_stage5[160]), .inData_161(wire_con_out_stage5[161]), .inData_162(wire_con_out_stage5[162]), .inData_163(wire_con_out_stage5[163]), .inData_164(wire_con_out_stage5[164]), .inData_165(wire_con_out_stage5[165]), .inData_166(wire_con_out_stage5[166]), .inData_167(wire_con_out_stage5[167]), .inData_168(wire_con_out_stage5[168]), .inData_169(wire_con_out_stage5[169]), .inData_170(wire_con_out_stage5[170]), .inData_171(wire_con_out_stage5[171]), .inData_172(wire_con_out_stage5[172]), .inData_173(wire_con_out_stage5[173]), .inData_174(wire_con_out_stage5[174]), .inData_175(wire_con_out_stage5[175]), .inData_176(wire_con_out_stage5[176]), .inData_177(wire_con_out_stage5[177]), .inData_178(wire_con_out_stage5[178]), .inData_179(wire_con_out_stage5[179]), .inData_180(wire_con_out_stage5[180]), .inData_181(wire_con_out_stage5[181]), .inData_182(wire_con_out_stage5[182]), .inData_183(wire_con_out_stage5[183]), .inData_184(wire_con_out_stage5[184]), .inData_185(wire_con_out_stage5[185]), .inData_186(wire_con_out_stage5[186]), .inData_187(wire_con_out_stage5[187]), .inData_188(wire_con_out_stage5[188]), .inData_189(wire_con_out_stage5[189]), .inData_190(wire_con_out_stage5[190]), .inData_191(wire_con_out_stage5[191]), .inData_192(wire_con_out_stage5[192]), .inData_193(wire_con_out_stage5[193]), .inData_194(wire_con_out_stage5[194]), .inData_195(wire_con_out_stage5[195]), .inData_196(wire_con_out_stage5[196]), .inData_197(wire_con_out_stage5[197]), .inData_198(wire_con_out_stage5[198]), .inData_199(wire_con_out_stage5[199]), .inData_200(wire_con_out_stage5[200]), .inData_201(wire_con_out_stage5[201]), .inData_202(wire_con_out_stage5[202]), .inData_203(wire_con_out_stage5[203]), .inData_204(wire_con_out_stage5[204]), .inData_205(wire_con_out_stage5[205]), .inData_206(wire_con_out_stage5[206]), .inData_207(wire_con_out_stage5[207]), .inData_208(wire_con_out_stage5[208]), .inData_209(wire_con_out_stage5[209]), .inData_210(wire_con_out_stage5[210]), .inData_211(wire_con_out_stage5[211]), .inData_212(wire_con_out_stage5[212]), .inData_213(wire_con_out_stage5[213]), .inData_214(wire_con_out_stage5[214]), .inData_215(wire_con_out_stage5[215]), .inData_216(wire_con_out_stage5[216]), .inData_217(wire_con_out_stage5[217]), .inData_218(wire_con_out_stage5[218]), .inData_219(wire_con_out_stage5[219]), .inData_220(wire_con_out_stage5[220]), .inData_221(wire_con_out_stage5[221]), .inData_222(wire_con_out_stage5[222]), .inData_223(wire_con_out_stage5[223]), .inData_224(wire_con_out_stage5[224]), .inData_225(wire_con_out_stage5[225]), .inData_226(wire_con_out_stage5[226]), .inData_227(wire_con_out_stage5[227]), .inData_228(wire_con_out_stage5[228]), .inData_229(wire_con_out_stage5[229]), .inData_230(wire_con_out_stage5[230]), .inData_231(wire_con_out_stage5[231]), .inData_232(wire_con_out_stage5[232]), .inData_233(wire_con_out_stage5[233]), .inData_234(wire_con_out_stage5[234]), .inData_235(wire_con_out_stage5[235]), .inData_236(wire_con_out_stage5[236]), .inData_237(wire_con_out_stage5[237]), .inData_238(wire_con_out_stage5[238]), .inData_239(wire_con_out_stage5[239]), .inData_240(wire_con_out_stage5[240]), .inData_241(wire_con_out_stage5[241]), .inData_242(wire_con_out_stage5[242]), .inData_243(wire_con_out_stage5[243]), .inData_244(wire_con_out_stage5[244]), .inData_245(wire_con_out_stage5[245]), .inData_246(wire_con_out_stage5[246]), .inData_247(wire_con_out_stage5[247]), .inData_248(wire_con_out_stage5[248]), .inData_249(wire_con_out_stage5[249]), .inData_250(wire_con_out_stage5[250]), .inData_251(wire_con_out_stage5[251]), .inData_252(wire_con_out_stage5[252]), .inData_253(wire_con_out_stage5[253]), .inData_254(wire_con_out_stage5[254]), .inData_255(wire_con_out_stage5[255]), 
        .outData_0(wire_con_in_stage6[0]), .outData_1(wire_con_in_stage6[1]), .outData_2(wire_con_in_stage6[2]), .outData_3(wire_con_in_stage6[3]), .outData_4(wire_con_in_stage6[4]), .outData_5(wire_con_in_stage6[5]), .outData_6(wire_con_in_stage6[6]), .outData_7(wire_con_in_stage6[7]), .outData_8(wire_con_in_stage6[8]), .outData_9(wire_con_in_stage6[9]), .outData_10(wire_con_in_stage6[10]), .outData_11(wire_con_in_stage6[11]), .outData_12(wire_con_in_stage6[12]), .outData_13(wire_con_in_stage6[13]), .outData_14(wire_con_in_stage6[14]), .outData_15(wire_con_in_stage6[15]), .outData_16(wire_con_in_stage6[16]), .outData_17(wire_con_in_stage6[17]), .outData_18(wire_con_in_stage6[18]), .outData_19(wire_con_in_stage6[19]), .outData_20(wire_con_in_stage6[20]), .outData_21(wire_con_in_stage6[21]), .outData_22(wire_con_in_stage6[22]), .outData_23(wire_con_in_stage6[23]), .outData_24(wire_con_in_stage6[24]), .outData_25(wire_con_in_stage6[25]), .outData_26(wire_con_in_stage6[26]), .outData_27(wire_con_in_stage6[27]), .outData_28(wire_con_in_stage6[28]), .outData_29(wire_con_in_stage6[29]), .outData_30(wire_con_in_stage6[30]), .outData_31(wire_con_in_stage6[31]), .outData_32(wire_con_in_stage6[32]), .outData_33(wire_con_in_stage6[33]), .outData_34(wire_con_in_stage6[34]), .outData_35(wire_con_in_stage6[35]), .outData_36(wire_con_in_stage6[36]), .outData_37(wire_con_in_stage6[37]), .outData_38(wire_con_in_stage6[38]), .outData_39(wire_con_in_stage6[39]), .outData_40(wire_con_in_stage6[40]), .outData_41(wire_con_in_stage6[41]), .outData_42(wire_con_in_stage6[42]), .outData_43(wire_con_in_stage6[43]), .outData_44(wire_con_in_stage6[44]), .outData_45(wire_con_in_stage6[45]), .outData_46(wire_con_in_stage6[46]), .outData_47(wire_con_in_stage6[47]), .outData_48(wire_con_in_stage6[48]), .outData_49(wire_con_in_stage6[49]), .outData_50(wire_con_in_stage6[50]), .outData_51(wire_con_in_stage6[51]), .outData_52(wire_con_in_stage6[52]), .outData_53(wire_con_in_stage6[53]), .outData_54(wire_con_in_stage6[54]), .outData_55(wire_con_in_stage6[55]), .outData_56(wire_con_in_stage6[56]), .outData_57(wire_con_in_stage6[57]), .outData_58(wire_con_in_stage6[58]), .outData_59(wire_con_in_stage6[59]), .outData_60(wire_con_in_stage6[60]), .outData_61(wire_con_in_stage6[61]), .outData_62(wire_con_in_stage6[62]), .outData_63(wire_con_in_stage6[63]), .outData_64(wire_con_in_stage6[64]), .outData_65(wire_con_in_stage6[65]), .outData_66(wire_con_in_stage6[66]), .outData_67(wire_con_in_stage6[67]), .outData_68(wire_con_in_stage6[68]), .outData_69(wire_con_in_stage6[69]), .outData_70(wire_con_in_stage6[70]), .outData_71(wire_con_in_stage6[71]), .outData_72(wire_con_in_stage6[72]), .outData_73(wire_con_in_stage6[73]), .outData_74(wire_con_in_stage6[74]), .outData_75(wire_con_in_stage6[75]), .outData_76(wire_con_in_stage6[76]), .outData_77(wire_con_in_stage6[77]), .outData_78(wire_con_in_stage6[78]), .outData_79(wire_con_in_stage6[79]), .outData_80(wire_con_in_stage6[80]), .outData_81(wire_con_in_stage6[81]), .outData_82(wire_con_in_stage6[82]), .outData_83(wire_con_in_stage6[83]), .outData_84(wire_con_in_stage6[84]), .outData_85(wire_con_in_stage6[85]), .outData_86(wire_con_in_stage6[86]), .outData_87(wire_con_in_stage6[87]), .outData_88(wire_con_in_stage6[88]), .outData_89(wire_con_in_stage6[89]), .outData_90(wire_con_in_stage6[90]), .outData_91(wire_con_in_stage6[91]), .outData_92(wire_con_in_stage6[92]), .outData_93(wire_con_in_stage6[93]), .outData_94(wire_con_in_stage6[94]), .outData_95(wire_con_in_stage6[95]), .outData_96(wire_con_in_stage6[96]), .outData_97(wire_con_in_stage6[97]), .outData_98(wire_con_in_stage6[98]), .outData_99(wire_con_in_stage6[99]), .outData_100(wire_con_in_stage6[100]), .outData_101(wire_con_in_stage6[101]), .outData_102(wire_con_in_stage6[102]), .outData_103(wire_con_in_stage6[103]), .outData_104(wire_con_in_stage6[104]), .outData_105(wire_con_in_stage6[105]), .outData_106(wire_con_in_stage6[106]), .outData_107(wire_con_in_stage6[107]), .outData_108(wire_con_in_stage6[108]), .outData_109(wire_con_in_stage6[109]), .outData_110(wire_con_in_stage6[110]), .outData_111(wire_con_in_stage6[111]), .outData_112(wire_con_in_stage6[112]), .outData_113(wire_con_in_stage6[113]), .outData_114(wire_con_in_stage6[114]), .outData_115(wire_con_in_stage6[115]), .outData_116(wire_con_in_stage6[116]), .outData_117(wire_con_in_stage6[117]), .outData_118(wire_con_in_stage6[118]), .outData_119(wire_con_in_stage6[119]), .outData_120(wire_con_in_stage6[120]), .outData_121(wire_con_in_stage6[121]), .outData_122(wire_con_in_stage6[122]), .outData_123(wire_con_in_stage6[123]), .outData_124(wire_con_in_stage6[124]), .outData_125(wire_con_in_stage6[125]), .outData_126(wire_con_in_stage6[126]), .outData_127(wire_con_in_stage6[127]), .outData_128(wire_con_in_stage6[128]), .outData_129(wire_con_in_stage6[129]), .outData_130(wire_con_in_stage6[130]), .outData_131(wire_con_in_stage6[131]), .outData_132(wire_con_in_stage6[132]), .outData_133(wire_con_in_stage6[133]), .outData_134(wire_con_in_stage6[134]), .outData_135(wire_con_in_stage6[135]), .outData_136(wire_con_in_stage6[136]), .outData_137(wire_con_in_stage6[137]), .outData_138(wire_con_in_stage6[138]), .outData_139(wire_con_in_stage6[139]), .outData_140(wire_con_in_stage6[140]), .outData_141(wire_con_in_stage6[141]), .outData_142(wire_con_in_stage6[142]), .outData_143(wire_con_in_stage6[143]), .outData_144(wire_con_in_stage6[144]), .outData_145(wire_con_in_stage6[145]), .outData_146(wire_con_in_stage6[146]), .outData_147(wire_con_in_stage6[147]), .outData_148(wire_con_in_stage6[148]), .outData_149(wire_con_in_stage6[149]), .outData_150(wire_con_in_stage6[150]), .outData_151(wire_con_in_stage6[151]), .outData_152(wire_con_in_stage6[152]), .outData_153(wire_con_in_stage6[153]), .outData_154(wire_con_in_stage6[154]), .outData_155(wire_con_in_stage6[155]), .outData_156(wire_con_in_stage6[156]), .outData_157(wire_con_in_stage6[157]), .outData_158(wire_con_in_stage6[158]), .outData_159(wire_con_in_stage6[159]), .outData_160(wire_con_in_stage6[160]), .outData_161(wire_con_in_stage6[161]), .outData_162(wire_con_in_stage6[162]), .outData_163(wire_con_in_stage6[163]), .outData_164(wire_con_in_stage6[164]), .outData_165(wire_con_in_stage6[165]), .outData_166(wire_con_in_stage6[166]), .outData_167(wire_con_in_stage6[167]), .outData_168(wire_con_in_stage6[168]), .outData_169(wire_con_in_stage6[169]), .outData_170(wire_con_in_stage6[170]), .outData_171(wire_con_in_stage6[171]), .outData_172(wire_con_in_stage6[172]), .outData_173(wire_con_in_stage6[173]), .outData_174(wire_con_in_stage6[174]), .outData_175(wire_con_in_stage6[175]), .outData_176(wire_con_in_stage6[176]), .outData_177(wire_con_in_stage6[177]), .outData_178(wire_con_in_stage6[178]), .outData_179(wire_con_in_stage6[179]), .outData_180(wire_con_in_stage6[180]), .outData_181(wire_con_in_stage6[181]), .outData_182(wire_con_in_stage6[182]), .outData_183(wire_con_in_stage6[183]), .outData_184(wire_con_in_stage6[184]), .outData_185(wire_con_in_stage6[185]), .outData_186(wire_con_in_stage6[186]), .outData_187(wire_con_in_stage6[187]), .outData_188(wire_con_in_stage6[188]), .outData_189(wire_con_in_stage6[189]), .outData_190(wire_con_in_stage6[190]), .outData_191(wire_con_in_stage6[191]), .outData_192(wire_con_in_stage6[192]), .outData_193(wire_con_in_stage6[193]), .outData_194(wire_con_in_stage6[194]), .outData_195(wire_con_in_stage6[195]), .outData_196(wire_con_in_stage6[196]), .outData_197(wire_con_in_stage6[197]), .outData_198(wire_con_in_stage6[198]), .outData_199(wire_con_in_stage6[199]), .outData_200(wire_con_in_stage6[200]), .outData_201(wire_con_in_stage6[201]), .outData_202(wire_con_in_stage6[202]), .outData_203(wire_con_in_stage6[203]), .outData_204(wire_con_in_stage6[204]), .outData_205(wire_con_in_stage6[205]), .outData_206(wire_con_in_stage6[206]), .outData_207(wire_con_in_stage6[207]), .outData_208(wire_con_in_stage6[208]), .outData_209(wire_con_in_stage6[209]), .outData_210(wire_con_in_stage6[210]), .outData_211(wire_con_in_stage6[211]), .outData_212(wire_con_in_stage6[212]), .outData_213(wire_con_in_stage6[213]), .outData_214(wire_con_in_stage6[214]), .outData_215(wire_con_in_stage6[215]), .outData_216(wire_con_in_stage6[216]), .outData_217(wire_con_in_stage6[217]), .outData_218(wire_con_in_stage6[218]), .outData_219(wire_con_in_stage6[219]), .outData_220(wire_con_in_stage6[220]), .outData_221(wire_con_in_stage6[221]), .outData_222(wire_con_in_stage6[222]), .outData_223(wire_con_in_stage6[223]), .outData_224(wire_con_in_stage6[224]), .outData_225(wire_con_in_stage6[225]), .outData_226(wire_con_in_stage6[226]), .outData_227(wire_con_in_stage6[227]), .outData_228(wire_con_in_stage6[228]), .outData_229(wire_con_in_stage6[229]), .outData_230(wire_con_in_stage6[230]), .outData_231(wire_con_in_stage6[231]), .outData_232(wire_con_in_stage6[232]), .outData_233(wire_con_in_stage6[233]), .outData_234(wire_con_in_stage6[234]), .outData_235(wire_con_in_stage6[235]), .outData_236(wire_con_in_stage6[236]), .outData_237(wire_con_in_stage6[237]), .outData_238(wire_con_in_stage6[238]), .outData_239(wire_con_in_stage6[239]), .outData_240(wire_con_in_stage6[240]), .outData_241(wire_con_in_stage6[241]), .outData_242(wire_con_in_stage6[242]), .outData_243(wire_con_in_stage6[243]), .outData_244(wire_con_in_stage6[244]), .outData_245(wire_con_in_stage6[245]), .outData_246(wire_con_in_stage6[246]), .outData_247(wire_con_in_stage6[247]), .outData_248(wire_con_in_stage6[248]), .outData_249(wire_con_in_stage6[249]), .outData_250(wire_con_in_stage6[250]), .outData_251(wire_con_in_stage6[251]), .outData_252(wire_con_in_stage6[252]), .outData_253(wire_con_in_stage6[253]), .outData_254(wire_con_in_stage6[254]), .outData_255(wire_con_in_stage6[255]), 
        .in_start(in_start_stage6), .out_start(con_in_start_stage6), .ctrl(wire_ctrl_stage6), .clk(clk), .rst(rst));
  
  wireCon_dp256_st6_L wire_stage_6(
        .inData_0(wire_con_in_stage6[0]), .inData_1(wire_con_in_stage6[1]), .inData_2(wire_con_in_stage6[2]), .inData_3(wire_con_in_stage6[3]), .inData_4(wire_con_in_stage6[4]), .inData_5(wire_con_in_stage6[5]), .inData_6(wire_con_in_stage6[6]), .inData_7(wire_con_in_stage6[7]), .inData_8(wire_con_in_stage6[8]), .inData_9(wire_con_in_stage6[9]), .inData_10(wire_con_in_stage6[10]), .inData_11(wire_con_in_stage6[11]), .inData_12(wire_con_in_stage6[12]), .inData_13(wire_con_in_stage6[13]), .inData_14(wire_con_in_stage6[14]), .inData_15(wire_con_in_stage6[15]), .inData_16(wire_con_in_stage6[16]), .inData_17(wire_con_in_stage6[17]), .inData_18(wire_con_in_stage6[18]), .inData_19(wire_con_in_stage6[19]), .inData_20(wire_con_in_stage6[20]), .inData_21(wire_con_in_stage6[21]), .inData_22(wire_con_in_stage6[22]), .inData_23(wire_con_in_stage6[23]), .inData_24(wire_con_in_stage6[24]), .inData_25(wire_con_in_stage6[25]), .inData_26(wire_con_in_stage6[26]), .inData_27(wire_con_in_stage6[27]), .inData_28(wire_con_in_stage6[28]), .inData_29(wire_con_in_stage6[29]), .inData_30(wire_con_in_stage6[30]), .inData_31(wire_con_in_stage6[31]), .inData_32(wire_con_in_stage6[32]), .inData_33(wire_con_in_stage6[33]), .inData_34(wire_con_in_stage6[34]), .inData_35(wire_con_in_stage6[35]), .inData_36(wire_con_in_stage6[36]), .inData_37(wire_con_in_stage6[37]), .inData_38(wire_con_in_stage6[38]), .inData_39(wire_con_in_stage6[39]), .inData_40(wire_con_in_stage6[40]), .inData_41(wire_con_in_stage6[41]), .inData_42(wire_con_in_stage6[42]), .inData_43(wire_con_in_stage6[43]), .inData_44(wire_con_in_stage6[44]), .inData_45(wire_con_in_stage6[45]), .inData_46(wire_con_in_stage6[46]), .inData_47(wire_con_in_stage6[47]), .inData_48(wire_con_in_stage6[48]), .inData_49(wire_con_in_stage6[49]), .inData_50(wire_con_in_stage6[50]), .inData_51(wire_con_in_stage6[51]), .inData_52(wire_con_in_stage6[52]), .inData_53(wire_con_in_stage6[53]), .inData_54(wire_con_in_stage6[54]), .inData_55(wire_con_in_stage6[55]), .inData_56(wire_con_in_stage6[56]), .inData_57(wire_con_in_stage6[57]), .inData_58(wire_con_in_stage6[58]), .inData_59(wire_con_in_stage6[59]), .inData_60(wire_con_in_stage6[60]), .inData_61(wire_con_in_stage6[61]), .inData_62(wire_con_in_stage6[62]), .inData_63(wire_con_in_stage6[63]), .inData_64(wire_con_in_stage6[64]), .inData_65(wire_con_in_stage6[65]), .inData_66(wire_con_in_stage6[66]), .inData_67(wire_con_in_stage6[67]), .inData_68(wire_con_in_stage6[68]), .inData_69(wire_con_in_stage6[69]), .inData_70(wire_con_in_stage6[70]), .inData_71(wire_con_in_stage6[71]), .inData_72(wire_con_in_stage6[72]), .inData_73(wire_con_in_stage6[73]), .inData_74(wire_con_in_stage6[74]), .inData_75(wire_con_in_stage6[75]), .inData_76(wire_con_in_stage6[76]), .inData_77(wire_con_in_stage6[77]), .inData_78(wire_con_in_stage6[78]), .inData_79(wire_con_in_stage6[79]), .inData_80(wire_con_in_stage6[80]), .inData_81(wire_con_in_stage6[81]), .inData_82(wire_con_in_stage6[82]), .inData_83(wire_con_in_stage6[83]), .inData_84(wire_con_in_stage6[84]), .inData_85(wire_con_in_stage6[85]), .inData_86(wire_con_in_stage6[86]), .inData_87(wire_con_in_stage6[87]), .inData_88(wire_con_in_stage6[88]), .inData_89(wire_con_in_stage6[89]), .inData_90(wire_con_in_stage6[90]), .inData_91(wire_con_in_stage6[91]), .inData_92(wire_con_in_stage6[92]), .inData_93(wire_con_in_stage6[93]), .inData_94(wire_con_in_stage6[94]), .inData_95(wire_con_in_stage6[95]), .inData_96(wire_con_in_stage6[96]), .inData_97(wire_con_in_stage6[97]), .inData_98(wire_con_in_stage6[98]), .inData_99(wire_con_in_stage6[99]), .inData_100(wire_con_in_stage6[100]), .inData_101(wire_con_in_stage6[101]), .inData_102(wire_con_in_stage6[102]), .inData_103(wire_con_in_stage6[103]), .inData_104(wire_con_in_stage6[104]), .inData_105(wire_con_in_stage6[105]), .inData_106(wire_con_in_stage6[106]), .inData_107(wire_con_in_stage6[107]), .inData_108(wire_con_in_stage6[108]), .inData_109(wire_con_in_stage6[109]), .inData_110(wire_con_in_stage6[110]), .inData_111(wire_con_in_stage6[111]), .inData_112(wire_con_in_stage6[112]), .inData_113(wire_con_in_stage6[113]), .inData_114(wire_con_in_stage6[114]), .inData_115(wire_con_in_stage6[115]), .inData_116(wire_con_in_stage6[116]), .inData_117(wire_con_in_stage6[117]), .inData_118(wire_con_in_stage6[118]), .inData_119(wire_con_in_stage6[119]), .inData_120(wire_con_in_stage6[120]), .inData_121(wire_con_in_stage6[121]), .inData_122(wire_con_in_stage6[122]), .inData_123(wire_con_in_stage6[123]), .inData_124(wire_con_in_stage6[124]), .inData_125(wire_con_in_stage6[125]), .inData_126(wire_con_in_stage6[126]), .inData_127(wire_con_in_stage6[127]), .inData_128(wire_con_in_stage6[128]), .inData_129(wire_con_in_stage6[129]), .inData_130(wire_con_in_stage6[130]), .inData_131(wire_con_in_stage6[131]), .inData_132(wire_con_in_stage6[132]), .inData_133(wire_con_in_stage6[133]), .inData_134(wire_con_in_stage6[134]), .inData_135(wire_con_in_stage6[135]), .inData_136(wire_con_in_stage6[136]), .inData_137(wire_con_in_stage6[137]), .inData_138(wire_con_in_stage6[138]), .inData_139(wire_con_in_stage6[139]), .inData_140(wire_con_in_stage6[140]), .inData_141(wire_con_in_stage6[141]), .inData_142(wire_con_in_stage6[142]), .inData_143(wire_con_in_stage6[143]), .inData_144(wire_con_in_stage6[144]), .inData_145(wire_con_in_stage6[145]), .inData_146(wire_con_in_stage6[146]), .inData_147(wire_con_in_stage6[147]), .inData_148(wire_con_in_stage6[148]), .inData_149(wire_con_in_stage6[149]), .inData_150(wire_con_in_stage6[150]), .inData_151(wire_con_in_stage6[151]), .inData_152(wire_con_in_stage6[152]), .inData_153(wire_con_in_stage6[153]), .inData_154(wire_con_in_stage6[154]), .inData_155(wire_con_in_stage6[155]), .inData_156(wire_con_in_stage6[156]), .inData_157(wire_con_in_stage6[157]), .inData_158(wire_con_in_stage6[158]), .inData_159(wire_con_in_stage6[159]), .inData_160(wire_con_in_stage6[160]), .inData_161(wire_con_in_stage6[161]), .inData_162(wire_con_in_stage6[162]), .inData_163(wire_con_in_stage6[163]), .inData_164(wire_con_in_stage6[164]), .inData_165(wire_con_in_stage6[165]), .inData_166(wire_con_in_stage6[166]), .inData_167(wire_con_in_stage6[167]), .inData_168(wire_con_in_stage6[168]), .inData_169(wire_con_in_stage6[169]), .inData_170(wire_con_in_stage6[170]), .inData_171(wire_con_in_stage6[171]), .inData_172(wire_con_in_stage6[172]), .inData_173(wire_con_in_stage6[173]), .inData_174(wire_con_in_stage6[174]), .inData_175(wire_con_in_stage6[175]), .inData_176(wire_con_in_stage6[176]), .inData_177(wire_con_in_stage6[177]), .inData_178(wire_con_in_stage6[178]), .inData_179(wire_con_in_stage6[179]), .inData_180(wire_con_in_stage6[180]), .inData_181(wire_con_in_stage6[181]), .inData_182(wire_con_in_stage6[182]), .inData_183(wire_con_in_stage6[183]), .inData_184(wire_con_in_stage6[184]), .inData_185(wire_con_in_stage6[185]), .inData_186(wire_con_in_stage6[186]), .inData_187(wire_con_in_stage6[187]), .inData_188(wire_con_in_stage6[188]), .inData_189(wire_con_in_stage6[189]), .inData_190(wire_con_in_stage6[190]), .inData_191(wire_con_in_stage6[191]), .inData_192(wire_con_in_stage6[192]), .inData_193(wire_con_in_stage6[193]), .inData_194(wire_con_in_stage6[194]), .inData_195(wire_con_in_stage6[195]), .inData_196(wire_con_in_stage6[196]), .inData_197(wire_con_in_stage6[197]), .inData_198(wire_con_in_stage6[198]), .inData_199(wire_con_in_stage6[199]), .inData_200(wire_con_in_stage6[200]), .inData_201(wire_con_in_stage6[201]), .inData_202(wire_con_in_stage6[202]), .inData_203(wire_con_in_stage6[203]), .inData_204(wire_con_in_stage6[204]), .inData_205(wire_con_in_stage6[205]), .inData_206(wire_con_in_stage6[206]), .inData_207(wire_con_in_stage6[207]), .inData_208(wire_con_in_stage6[208]), .inData_209(wire_con_in_stage6[209]), .inData_210(wire_con_in_stage6[210]), .inData_211(wire_con_in_stage6[211]), .inData_212(wire_con_in_stage6[212]), .inData_213(wire_con_in_stage6[213]), .inData_214(wire_con_in_stage6[214]), .inData_215(wire_con_in_stage6[215]), .inData_216(wire_con_in_stage6[216]), .inData_217(wire_con_in_stage6[217]), .inData_218(wire_con_in_stage6[218]), .inData_219(wire_con_in_stage6[219]), .inData_220(wire_con_in_stage6[220]), .inData_221(wire_con_in_stage6[221]), .inData_222(wire_con_in_stage6[222]), .inData_223(wire_con_in_stage6[223]), .inData_224(wire_con_in_stage6[224]), .inData_225(wire_con_in_stage6[225]), .inData_226(wire_con_in_stage6[226]), .inData_227(wire_con_in_stage6[227]), .inData_228(wire_con_in_stage6[228]), .inData_229(wire_con_in_stage6[229]), .inData_230(wire_con_in_stage6[230]), .inData_231(wire_con_in_stage6[231]), .inData_232(wire_con_in_stage6[232]), .inData_233(wire_con_in_stage6[233]), .inData_234(wire_con_in_stage6[234]), .inData_235(wire_con_in_stage6[235]), .inData_236(wire_con_in_stage6[236]), .inData_237(wire_con_in_stage6[237]), .inData_238(wire_con_in_stage6[238]), .inData_239(wire_con_in_stage6[239]), .inData_240(wire_con_in_stage6[240]), .inData_241(wire_con_in_stage6[241]), .inData_242(wire_con_in_stage6[242]), .inData_243(wire_con_in_stage6[243]), .inData_244(wire_con_in_stage6[244]), .inData_245(wire_con_in_stage6[245]), .inData_246(wire_con_in_stage6[246]), .inData_247(wire_con_in_stage6[247]), .inData_248(wire_con_in_stage6[248]), .inData_249(wire_con_in_stage6[249]), .inData_250(wire_con_in_stage6[250]), .inData_251(wire_con_in_stage6[251]), .inData_252(wire_con_in_stage6[252]), .inData_253(wire_con_in_stage6[253]), .inData_254(wire_con_in_stage6[254]), .inData_255(wire_con_in_stage6[255]), 
        .outData_0(wire_con_out_stage6[0]), .outData_1(wire_con_out_stage6[1]), .outData_2(wire_con_out_stage6[2]), .outData_3(wire_con_out_stage6[3]), .outData_4(wire_con_out_stage6[4]), .outData_5(wire_con_out_stage6[5]), .outData_6(wire_con_out_stage6[6]), .outData_7(wire_con_out_stage6[7]), .outData_8(wire_con_out_stage6[8]), .outData_9(wire_con_out_stage6[9]), .outData_10(wire_con_out_stage6[10]), .outData_11(wire_con_out_stage6[11]), .outData_12(wire_con_out_stage6[12]), .outData_13(wire_con_out_stage6[13]), .outData_14(wire_con_out_stage6[14]), .outData_15(wire_con_out_stage6[15]), .outData_16(wire_con_out_stage6[16]), .outData_17(wire_con_out_stage6[17]), .outData_18(wire_con_out_stage6[18]), .outData_19(wire_con_out_stage6[19]), .outData_20(wire_con_out_stage6[20]), .outData_21(wire_con_out_stage6[21]), .outData_22(wire_con_out_stage6[22]), .outData_23(wire_con_out_stage6[23]), .outData_24(wire_con_out_stage6[24]), .outData_25(wire_con_out_stage6[25]), .outData_26(wire_con_out_stage6[26]), .outData_27(wire_con_out_stage6[27]), .outData_28(wire_con_out_stage6[28]), .outData_29(wire_con_out_stage6[29]), .outData_30(wire_con_out_stage6[30]), .outData_31(wire_con_out_stage6[31]), .outData_32(wire_con_out_stage6[32]), .outData_33(wire_con_out_stage6[33]), .outData_34(wire_con_out_stage6[34]), .outData_35(wire_con_out_stage6[35]), .outData_36(wire_con_out_stage6[36]), .outData_37(wire_con_out_stage6[37]), .outData_38(wire_con_out_stage6[38]), .outData_39(wire_con_out_stage6[39]), .outData_40(wire_con_out_stage6[40]), .outData_41(wire_con_out_stage6[41]), .outData_42(wire_con_out_stage6[42]), .outData_43(wire_con_out_stage6[43]), .outData_44(wire_con_out_stage6[44]), .outData_45(wire_con_out_stage6[45]), .outData_46(wire_con_out_stage6[46]), .outData_47(wire_con_out_stage6[47]), .outData_48(wire_con_out_stage6[48]), .outData_49(wire_con_out_stage6[49]), .outData_50(wire_con_out_stage6[50]), .outData_51(wire_con_out_stage6[51]), .outData_52(wire_con_out_stage6[52]), .outData_53(wire_con_out_stage6[53]), .outData_54(wire_con_out_stage6[54]), .outData_55(wire_con_out_stage6[55]), .outData_56(wire_con_out_stage6[56]), .outData_57(wire_con_out_stage6[57]), .outData_58(wire_con_out_stage6[58]), .outData_59(wire_con_out_stage6[59]), .outData_60(wire_con_out_stage6[60]), .outData_61(wire_con_out_stage6[61]), .outData_62(wire_con_out_stage6[62]), .outData_63(wire_con_out_stage6[63]), .outData_64(wire_con_out_stage6[64]), .outData_65(wire_con_out_stage6[65]), .outData_66(wire_con_out_stage6[66]), .outData_67(wire_con_out_stage6[67]), .outData_68(wire_con_out_stage6[68]), .outData_69(wire_con_out_stage6[69]), .outData_70(wire_con_out_stage6[70]), .outData_71(wire_con_out_stage6[71]), .outData_72(wire_con_out_stage6[72]), .outData_73(wire_con_out_stage6[73]), .outData_74(wire_con_out_stage6[74]), .outData_75(wire_con_out_stage6[75]), .outData_76(wire_con_out_stage6[76]), .outData_77(wire_con_out_stage6[77]), .outData_78(wire_con_out_stage6[78]), .outData_79(wire_con_out_stage6[79]), .outData_80(wire_con_out_stage6[80]), .outData_81(wire_con_out_stage6[81]), .outData_82(wire_con_out_stage6[82]), .outData_83(wire_con_out_stage6[83]), .outData_84(wire_con_out_stage6[84]), .outData_85(wire_con_out_stage6[85]), .outData_86(wire_con_out_stage6[86]), .outData_87(wire_con_out_stage6[87]), .outData_88(wire_con_out_stage6[88]), .outData_89(wire_con_out_stage6[89]), .outData_90(wire_con_out_stage6[90]), .outData_91(wire_con_out_stage6[91]), .outData_92(wire_con_out_stage6[92]), .outData_93(wire_con_out_stage6[93]), .outData_94(wire_con_out_stage6[94]), .outData_95(wire_con_out_stage6[95]), .outData_96(wire_con_out_stage6[96]), .outData_97(wire_con_out_stage6[97]), .outData_98(wire_con_out_stage6[98]), .outData_99(wire_con_out_stage6[99]), .outData_100(wire_con_out_stage6[100]), .outData_101(wire_con_out_stage6[101]), .outData_102(wire_con_out_stage6[102]), .outData_103(wire_con_out_stage6[103]), .outData_104(wire_con_out_stage6[104]), .outData_105(wire_con_out_stage6[105]), .outData_106(wire_con_out_stage6[106]), .outData_107(wire_con_out_stage6[107]), .outData_108(wire_con_out_stage6[108]), .outData_109(wire_con_out_stage6[109]), .outData_110(wire_con_out_stage6[110]), .outData_111(wire_con_out_stage6[111]), .outData_112(wire_con_out_stage6[112]), .outData_113(wire_con_out_stage6[113]), .outData_114(wire_con_out_stage6[114]), .outData_115(wire_con_out_stage6[115]), .outData_116(wire_con_out_stage6[116]), .outData_117(wire_con_out_stage6[117]), .outData_118(wire_con_out_stage6[118]), .outData_119(wire_con_out_stage6[119]), .outData_120(wire_con_out_stage6[120]), .outData_121(wire_con_out_stage6[121]), .outData_122(wire_con_out_stage6[122]), .outData_123(wire_con_out_stage6[123]), .outData_124(wire_con_out_stage6[124]), .outData_125(wire_con_out_stage6[125]), .outData_126(wire_con_out_stage6[126]), .outData_127(wire_con_out_stage6[127]), .outData_128(wire_con_out_stage6[128]), .outData_129(wire_con_out_stage6[129]), .outData_130(wire_con_out_stage6[130]), .outData_131(wire_con_out_stage6[131]), .outData_132(wire_con_out_stage6[132]), .outData_133(wire_con_out_stage6[133]), .outData_134(wire_con_out_stage6[134]), .outData_135(wire_con_out_stage6[135]), .outData_136(wire_con_out_stage6[136]), .outData_137(wire_con_out_stage6[137]), .outData_138(wire_con_out_stage6[138]), .outData_139(wire_con_out_stage6[139]), .outData_140(wire_con_out_stage6[140]), .outData_141(wire_con_out_stage6[141]), .outData_142(wire_con_out_stage6[142]), .outData_143(wire_con_out_stage6[143]), .outData_144(wire_con_out_stage6[144]), .outData_145(wire_con_out_stage6[145]), .outData_146(wire_con_out_stage6[146]), .outData_147(wire_con_out_stage6[147]), .outData_148(wire_con_out_stage6[148]), .outData_149(wire_con_out_stage6[149]), .outData_150(wire_con_out_stage6[150]), .outData_151(wire_con_out_stage6[151]), .outData_152(wire_con_out_stage6[152]), .outData_153(wire_con_out_stage6[153]), .outData_154(wire_con_out_stage6[154]), .outData_155(wire_con_out_stage6[155]), .outData_156(wire_con_out_stage6[156]), .outData_157(wire_con_out_stage6[157]), .outData_158(wire_con_out_stage6[158]), .outData_159(wire_con_out_stage6[159]), .outData_160(wire_con_out_stage6[160]), .outData_161(wire_con_out_stage6[161]), .outData_162(wire_con_out_stage6[162]), .outData_163(wire_con_out_stage6[163]), .outData_164(wire_con_out_stage6[164]), .outData_165(wire_con_out_stage6[165]), .outData_166(wire_con_out_stage6[166]), .outData_167(wire_con_out_stage6[167]), .outData_168(wire_con_out_stage6[168]), .outData_169(wire_con_out_stage6[169]), .outData_170(wire_con_out_stage6[170]), .outData_171(wire_con_out_stage6[171]), .outData_172(wire_con_out_stage6[172]), .outData_173(wire_con_out_stage6[173]), .outData_174(wire_con_out_stage6[174]), .outData_175(wire_con_out_stage6[175]), .outData_176(wire_con_out_stage6[176]), .outData_177(wire_con_out_stage6[177]), .outData_178(wire_con_out_stage6[178]), .outData_179(wire_con_out_stage6[179]), .outData_180(wire_con_out_stage6[180]), .outData_181(wire_con_out_stage6[181]), .outData_182(wire_con_out_stage6[182]), .outData_183(wire_con_out_stage6[183]), .outData_184(wire_con_out_stage6[184]), .outData_185(wire_con_out_stage6[185]), .outData_186(wire_con_out_stage6[186]), .outData_187(wire_con_out_stage6[187]), .outData_188(wire_con_out_stage6[188]), .outData_189(wire_con_out_stage6[189]), .outData_190(wire_con_out_stage6[190]), .outData_191(wire_con_out_stage6[191]), .outData_192(wire_con_out_stage6[192]), .outData_193(wire_con_out_stage6[193]), .outData_194(wire_con_out_stage6[194]), .outData_195(wire_con_out_stage6[195]), .outData_196(wire_con_out_stage6[196]), .outData_197(wire_con_out_stage6[197]), .outData_198(wire_con_out_stage6[198]), .outData_199(wire_con_out_stage6[199]), .outData_200(wire_con_out_stage6[200]), .outData_201(wire_con_out_stage6[201]), .outData_202(wire_con_out_stage6[202]), .outData_203(wire_con_out_stage6[203]), .outData_204(wire_con_out_stage6[204]), .outData_205(wire_con_out_stage6[205]), .outData_206(wire_con_out_stage6[206]), .outData_207(wire_con_out_stage6[207]), .outData_208(wire_con_out_stage6[208]), .outData_209(wire_con_out_stage6[209]), .outData_210(wire_con_out_stage6[210]), .outData_211(wire_con_out_stage6[211]), .outData_212(wire_con_out_stage6[212]), .outData_213(wire_con_out_stage6[213]), .outData_214(wire_con_out_stage6[214]), .outData_215(wire_con_out_stage6[215]), .outData_216(wire_con_out_stage6[216]), .outData_217(wire_con_out_stage6[217]), .outData_218(wire_con_out_stage6[218]), .outData_219(wire_con_out_stage6[219]), .outData_220(wire_con_out_stage6[220]), .outData_221(wire_con_out_stage6[221]), .outData_222(wire_con_out_stage6[222]), .outData_223(wire_con_out_stage6[223]), .outData_224(wire_con_out_stage6[224]), .outData_225(wire_con_out_stage6[225]), .outData_226(wire_con_out_stage6[226]), .outData_227(wire_con_out_stage6[227]), .outData_228(wire_con_out_stage6[228]), .outData_229(wire_con_out_stage6[229]), .outData_230(wire_con_out_stage6[230]), .outData_231(wire_con_out_stage6[231]), .outData_232(wire_con_out_stage6[232]), .outData_233(wire_con_out_stage6[233]), .outData_234(wire_con_out_stage6[234]), .outData_235(wire_con_out_stage6[235]), .outData_236(wire_con_out_stage6[236]), .outData_237(wire_con_out_stage6[237]), .outData_238(wire_con_out_stage6[238]), .outData_239(wire_con_out_stage6[239]), .outData_240(wire_con_out_stage6[240]), .outData_241(wire_con_out_stage6[241]), .outData_242(wire_con_out_stage6[242]), .outData_243(wire_con_out_stage6[243]), .outData_244(wire_con_out_stage6[244]), .outData_245(wire_con_out_stage6[245]), .outData_246(wire_con_out_stage6[246]), .outData_247(wire_con_out_stage6[247]), .outData_248(wire_con_out_stage6[248]), .outData_249(wire_con_out_stage6[249]), .outData_250(wire_con_out_stage6[250]), .outData_251(wire_con_out_stage6[251]), .outData_252(wire_con_out_stage6[252]), .outData_253(wire_con_out_stage6[253]), .outData_254(wire_con_out_stage6[254]), .outData_255(wire_con_out_stage6[255]), 
        .in_start(con_in_start_stage6), .out_start(in_start_stage7), .clk(clk), .rst(rst)); 

  
  assign wire_ctrl_stage6[0] = counter_w[1]; 
  assign wire_ctrl_stage6[1] = counter_w[1]; 
  assign wire_ctrl_stage6[2] = counter_w[1]; 
  assign wire_ctrl_stage6[3] = counter_w[1]; 
  assign wire_ctrl_stage6[4] = counter_w[1]; 
  assign wire_ctrl_stage6[5] = counter_w[1]; 
  assign wire_ctrl_stage6[6] = counter_w[1]; 
  assign wire_ctrl_stage6[7] = counter_w[1]; 
  assign wire_ctrl_stage6[8] = counter_w[1]; 
  assign wire_ctrl_stage6[9] = counter_w[1]; 
  assign wire_ctrl_stage6[10] = counter_w[1]; 
  assign wire_ctrl_stage6[11] = counter_w[1]; 
  assign wire_ctrl_stage6[12] = counter_w[1]; 
  assign wire_ctrl_stage6[13] = counter_w[1]; 
  assign wire_ctrl_stage6[14] = counter_w[1]; 
  assign wire_ctrl_stage6[15] = counter_w[1]; 
  assign wire_ctrl_stage6[16] = counter_w[1]; 
  assign wire_ctrl_stage6[17] = counter_w[1]; 
  assign wire_ctrl_stage6[18] = counter_w[1]; 
  assign wire_ctrl_stage6[19] = counter_w[1]; 
  assign wire_ctrl_stage6[20] = counter_w[1]; 
  assign wire_ctrl_stage6[21] = counter_w[1]; 
  assign wire_ctrl_stage6[22] = counter_w[1]; 
  assign wire_ctrl_stage6[23] = counter_w[1]; 
  assign wire_ctrl_stage6[24] = counter_w[1]; 
  assign wire_ctrl_stage6[25] = counter_w[1]; 
  assign wire_ctrl_stage6[26] = counter_w[1]; 
  assign wire_ctrl_stage6[27] = counter_w[1]; 
  assign wire_ctrl_stage6[28] = counter_w[1]; 
  assign wire_ctrl_stage6[29] = counter_w[1]; 
  assign wire_ctrl_stage6[30] = counter_w[1]; 
  assign wire_ctrl_stage6[31] = counter_w[1]; 
  assign wire_ctrl_stage6[32] = counter_w[1]; 
  assign wire_ctrl_stage6[33] = counter_w[1]; 
  assign wire_ctrl_stage6[34] = counter_w[1]; 
  assign wire_ctrl_stage6[35] = counter_w[1]; 
  assign wire_ctrl_stage6[36] = counter_w[1]; 
  assign wire_ctrl_stage6[37] = counter_w[1]; 
  assign wire_ctrl_stage6[38] = counter_w[1]; 
  assign wire_ctrl_stage6[39] = counter_w[1]; 
  assign wire_ctrl_stage6[40] = counter_w[1]; 
  assign wire_ctrl_stage6[41] = counter_w[1]; 
  assign wire_ctrl_stage6[42] = counter_w[1]; 
  assign wire_ctrl_stage6[43] = counter_w[1]; 
  assign wire_ctrl_stage6[44] = counter_w[1]; 
  assign wire_ctrl_stage6[45] = counter_w[1]; 
  assign wire_ctrl_stage6[46] = counter_w[1]; 
  assign wire_ctrl_stage6[47] = counter_w[1]; 
  assign wire_ctrl_stage6[48] = counter_w[1]; 
  assign wire_ctrl_stage6[49] = counter_w[1]; 
  assign wire_ctrl_stage6[50] = counter_w[1]; 
  assign wire_ctrl_stage6[51] = counter_w[1]; 
  assign wire_ctrl_stage6[52] = counter_w[1]; 
  assign wire_ctrl_stage6[53] = counter_w[1]; 
  assign wire_ctrl_stage6[54] = counter_w[1]; 
  assign wire_ctrl_stage6[55] = counter_w[1]; 
  assign wire_ctrl_stage6[56] = counter_w[1]; 
  assign wire_ctrl_stage6[57] = counter_w[1]; 
  assign wire_ctrl_stage6[58] = counter_w[1]; 
  assign wire_ctrl_stage6[59] = counter_w[1]; 
  assign wire_ctrl_stage6[60] = counter_w[1]; 
  assign wire_ctrl_stage6[61] = counter_w[1]; 
  assign wire_ctrl_stage6[62] = counter_w[1]; 
  assign wire_ctrl_stage6[63] = counter_w[1]; 
  assign wire_ctrl_stage6[64] = counter_w[1]; 
  assign wire_ctrl_stage6[65] = counter_w[1]; 
  assign wire_ctrl_stage6[66] = counter_w[1]; 
  assign wire_ctrl_stage6[67] = counter_w[1]; 
  assign wire_ctrl_stage6[68] = counter_w[1]; 
  assign wire_ctrl_stage6[69] = counter_w[1]; 
  assign wire_ctrl_stage6[70] = counter_w[1]; 
  assign wire_ctrl_stage6[71] = counter_w[1]; 
  assign wire_ctrl_stage6[72] = counter_w[1]; 
  assign wire_ctrl_stage6[73] = counter_w[1]; 
  assign wire_ctrl_stage6[74] = counter_w[1]; 
  assign wire_ctrl_stage6[75] = counter_w[1]; 
  assign wire_ctrl_stage6[76] = counter_w[1]; 
  assign wire_ctrl_stage6[77] = counter_w[1]; 
  assign wire_ctrl_stage6[78] = counter_w[1]; 
  assign wire_ctrl_stage6[79] = counter_w[1]; 
  assign wire_ctrl_stage6[80] = counter_w[1]; 
  assign wire_ctrl_stage6[81] = counter_w[1]; 
  assign wire_ctrl_stage6[82] = counter_w[1]; 
  assign wire_ctrl_stage6[83] = counter_w[1]; 
  assign wire_ctrl_stage6[84] = counter_w[1]; 
  assign wire_ctrl_stage6[85] = counter_w[1]; 
  assign wire_ctrl_stage6[86] = counter_w[1]; 
  assign wire_ctrl_stage6[87] = counter_w[1]; 
  assign wire_ctrl_stage6[88] = counter_w[1]; 
  assign wire_ctrl_stage6[89] = counter_w[1]; 
  assign wire_ctrl_stage6[90] = counter_w[1]; 
  assign wire_ctrl_stage6[91] = counter_w[1]; 
  assign wire_ctrl_stage6[92] = counter_w[1]; 
  assign wire_ctrl_stage6[93] = counter_w[1]; 
  assign wire_ctrl_stage6[94] = counter_w[1]; 
  assign wire_ctrl_stage6[95] = counter_w[1]; 
  assign wire_ctrl_stage6[96] = counter_w[1]; 
  assign wire_ctrl_stage6[97] = counter_w[1]; 
  assign wire_ctrl_stage6[98] = counter_w[1]; 
  assign wire_ctrl_stage6[99] = counter_w[1]; 
  assign wire_ctrl_stage6[100] = counter_w[1]; 
  assign wire_ctrl_stage6[101] = counter_w[1]; 
  assign wire_ctrl_stage6[102] = counter_w[1]; 
  assign wire_ctrl_stage6[103] = counter_w[1]; 
  assign wire_ctrl_stage6[104] = counter_w[1]; 
  assign wire_ctrl_stage6[105] = counter_w[1]; 
  assign wire_ctrl_stage6[106] = counter_w[1]; 
  assign wire_ctrl_stage6[107] = counter_w[1]; 
  assign wire_ctrl_stage6[108] = counter_w[1]; 
  assign wire_ctrl_stage6[109] = counter_w[1]; 
  assign wire_ctrl_stage6[110] = counter_w[1]; 
  assign wire_ctrl_stage6[111] = counter_w[1]; 
  assign wire_ctrl_stage6[112] = counter_w[1]; 
  assign wire_ctrl_stage6[113] = counter_w[1]; 
  assign wire_ctrl_stage6[114] = counter_w[1]; 
  assign wire_ctrl_stage6[115] = counter_w[1]; 
  assign wire_ctrl_stage6[116] = counter_w[1]; 
  assign wire_ctrl_stage6[117] = counter_w[1]; 
  assign wire_ctrl_stage6[118] = counter_w[1]; 
  assign wire_ctrl_stage6[119] = counter_w[1]; 
  assign wire_ctrl_stage6[120] = counter_w[1]; 
  assign wire_ctrl_stage6[121] = counter_w[1]; 
  assign wire_ctrl_stage6[122] = counter_w[1]; 
  assign wire_ctrl_stage6[123] = counter_w[1]; 
  assign wire_ctrl_stage6[124] = counter_w[1]; 
  assign wire_ctrl_stage6[125] = counter_w[1]; 
  assign wire_ctrl_stage6[126] = counter_w[1]; 
  assign wire_ctrl_stage6[127] = counter_w[1]; 
  wire [DATA_WIDTH-1:0] wire_con_in_stage7[255:0];
  wire [DATA_WIDTH-1:0] wire_con_out_stage7[255:0];
  wire [127:0] wire_ctrl_stage7;

  switches_stage_st7_0_L switch_stage_7(
        .inData_0(wire_con_out_stage6[0]), .inData_1(wire_con_out_stage6[1]), .inData_2(wire_con_out_stage6[2]), .inData_3(wire_con_out_stage6[3]), .inData_4(wire_con_out_stage6[4]), .inData_5(wire_con_out_stage6[5]), .inData_6(wire_con_out_stage6[6]), .inData_7(wire_con_out_stage6[7]), .inData_8(wire_con_out_stage6[8]), .inData_9(wire_con_out_stage6[9]), .inData_10(wire_con_out_stage6[10]), .inData_11(wire_con_out_stage6[11]), .inData_12(wire_con_out_stage6[12]), .inData_13(wire_con_out_stage6[13]), .inData_14(wire_con_out_stage6[14]), .inData_15(wire_con_out_stage6[15]), .inData_16(wire_con_out_stage6[16]), .inData_17(wire_con_out_stage6[17]), .inData_18(wire_con_out_stage6[18]), .inData_19(wire_con_out_stage6[19]), .inData_20(wire_con_out_stage6[20]), .inData_21(wire_con_out_stage6[21]), .inData_22(wire_con_out_stage6[22]), .inData_23(wire_con_out_stage6[23]), .inData_24(wire_con_out_stage6[24]), .inData_25(wire_con_out_stage6[25]), .inData_26(wire_con_out_stage6[26]), .inData_27(wire_con_out_stage6[27]), .inData_28(wire_con_out_stage6[28]), .inData_29(wire_con_out_stage6[29]), .inData_30(wire_con_out_stage6[30]), .inData_31(wire_con_out_stage6[31]), .inData_32(wire_con_out_stage6[32]), .inData_33(wire_con_out_stage6[33]), .inData_34(wire_con_out_stage6[34]), .inData_35(wire_con_out_stage6[35]), .inData_36(wire_con_out_stage6[36]), .inData_37(wire_con_out_stage6[37]), .inData_38(wire_con_out_stage6[38]), .inData_39(wire_con_out_stage6[39]), .inData_40(wire_con_out_stage6[40]), .inData_41(wire_con_out_stage6[41]), .inData_42(wire_con_out_stage6[42]), .inData_43(wire_con_out_stage6[43]), .inData_44(wire_con_out_stage6[44]), .inData_45(wire_con_out_stage6[45]), .inData_46(wire_con_out_stage6[46]), .inData_47(wire_con_out_stage6[47]), .inData_48(wire_con_out_stage6[48]), .inData_49(wire_con_out_stage6[49]), .inData_50(wire_con_out_stage6[50]), .inData_51(wire_con_out_stage6[51]), .inData_52(wire_con_out_stage6[52]), .inData_53(wire_con_out_stage6[53]), .inData_54(wire_con_out_stage6[54]), .inData_55(wire_con_out_stage6[55]), .inData_56(wire_con_out_stage6[56]), .inData_57(wire_con_out_stage6[57]), .inData_58(wire_con_out_stage6[58]), .inData_59(wire_con_out_stage6[59]), .inData_60(wire_con_out_stage6[60]), .inData_61(wire_con_out_stage6[61]), .inData_62(wire_con_out_stage6[62]), .inData_63(wire_con_out_stage6[63]), .inData_64(wire_con_out_stage6[64]), .inData_65(wire_con_out_stage6[65]), .inData_66(wire_con_out_stage6[66]), .inData_67(wire_con_out_stage6[67]), .inData_68(wire_con_out_stage6[68]), .inData_69(wire_con_out_stage6[69]), .inData_70(wire_con_out_stage6[70]), .inData_71(wire_con_out_stage6[71]), .inData_72(wire_con_out_stage6[72]), .inData_73(wire_con_out_stage6[73]), .inData_74(wire_con_out_stage6[74]), .inData_75(wire_con_out_stage6[75]), .inData_76(wire_con_out_stage6[76]), .inData_77(wire_con_out_stage6[77]), .inData_78(wire_con_out_stage6[78]), .inData_79(wire_con_out_stage6[79]), .inData_80(wire_con_out_stage6[80]), .inData_81(wire_con_out_stage6[81]), .inData_82(wire_con_out_stage6[82]), .inData_83(wire_con_out_stage6[83]), .inData_84(wire_con_out_stage6[84]), .inData_85(wire_con_out_stage6[85]), .inData_86(wire_con_out_stage6[86]), .inData_87(wire_con_out_stage6[87]), .inData_88(wire_con_out_stage6[88]), .inData_89(wire_con_out_stage6[89]), .inData_90(wire_con_out_stage6[90]), .inData_91(wire_con_out_stage6[91]), .inData_92(wire_con_out_stage6[92]), .inData_93(wire_con_out_stage6[93]), .inData_94(wire_con_out_stage6[94]), .inData_95(wire_con_out_stage6[95]), .inData_96(wire_con_out_stage6[96]), .inData_97(wire_con_out_stage6[97]), .inData_98(wire_con_out_stage6[98]), .inData_99(wire_con_out_stage6[99]), .inData_100(wire_con_out_stage6[100]), .inData_101(wire_con_out_stage6[101]), .inData_102(wire_con_out_stage6[102]), .inData_103(wire_con_out_stage6[103]), .inData_104(wire_con_out_stage6[104]), .inData_105(wire_con_out_stage6[105]), .inData_106(wire_con_out_stage6[106]), .inData_107(wire_con_out_stage6[107]), .inData_108(wire_con_out_stage6[108]), .inData_109(wire_con_out_stage6[109]), .inData_110(wire_con_out_stage6[110]), .inData_111(wire_con_out_stage6[111]), .inData_112(wire_con_out_stage6[112]), .inData_113(wire_con_out_stage6[113]), .inData_114(wire_con_out_stage6[114]), .inData_115(wire_con_out_stage6[115]), .inData_116(wire_con_out_stage6[116]), .inData_117(wire_con_out_stage6[117]), .inData_118(wire_con_out_stage6[118]), .inData_119(wire_con_out_stage6[119]), .inData_120(wire_con_out_stage6[120]), .inData_121(wire_con_out_stage6[121]), .inData_122(wire_con_out_stage6[122]), .inData_123(wire_con_out_stage6[123]), .inData_124(wire_con_out_stage6[124]), .inData_125(wire_con_out_stage6[125]), .inData_126(wire_con_out_stage6[126]), .inData_127(wire_con_out_stage6[127]), .inData_128(wire_con_out_stage6[128]), .inData_129(wire_con_out_stage6[129]), .inData_130(wire_con_out_stage6[130]), .inData_131(wire_con_out_stage6[131]), .inData_132(wire_con_out_stage6[132]), .inData_133(wire_con_out_stage6[133]), .inData_134(wire_con_out_stage6[134]), .inData_135(wire_con_out_stage6[135]), .inData_136(wire_con_out_stage6[136]), .inData_137(wire_con_out_stage6[137]), .inData_138(wire_con_out_stage6[138]), .inData_139(wire_con_out_stage6[139]), .inData_140(wire_con_out_stage6[140]), .inData_141(wire_con_out_stage6[141]), .inData_142(wire_con_out_stage6[142]), .inData_143(wire_con_out_stage6[143]), .inData_144(wire_con_out_stage6[144]), .inData_145(wire_con_out_stage6[145]), .inData_146(wire_con_out_stage6[146]), .inData_147(wire_con_out_stage6[147]), .inData_148(wire_con_out_stage6[148]), .inData_149(wire_con_out_stage6[149]), .inData_150(wire_con_out_stage6[150]), .inData_151(wire_con_out_stage6[151]), .inData_152(wire_con_out_stage6[152]), .inData_153(wire_con_out_stage6[153]), .inData_154(wire_con_out_stage6[154]), .inData_155(wire_con_out_stage6[155]), .inData_156(wire_con_out_stage6[156]), .inData_157(wire_con_out_stage6[157]), .inData_158(wire_con_out_stage6[158]), .inData_159(wire_con_out_stage6[159]), .inData_160(wire_con_out_stage6[160]), .inData_161(wire_con_out_stage6[161]), .inData_162(wire_con_out_stage6[162]), .inData_163(wire_con_out_stage6[163]), .inData_164(wire_con_out_stage6[164]), .inData_165(wire_con_out_stage6[165]), .inData_166(wire_con_out_stage6[166]), .inData_167(wire_con_out_stage6[167]), .inData_168(wire_con_out_stage6[168]), .inData_169(wire_con_out_stage6[169]), .inData_170(wire_con_out_stage6[170]), .inData_171(wire_con_out_stage6[171]), .inData_172(wire_con_out_stage6[172]), .inData_173(wire_con_out_stage6[173]), .inData_174(wire_con_out_stage6[174]), .inData_175(wire_con_out_stage6[175]), .inData_176(wire_con_out_stage6[176]), .inData_177(wire_con_out_stage6[177]), .inData_178(wire_con_out_stage6[178]), .inData_179(wire_con_out_stage6[179]), .inData_180(wire_con_out_stage6[180]), .inData_181(wire_con_out_stage6[181]), .inData_182(wire_con_out_stage6[182]), .inData_183(wire_con_out_stage6[183]), .inData_184(wire_con_out_stage6[184]), .inData_185(wire_con_out_stage6[185]), .inData_186(wire_con_out_stage6[186]), .inData_187(wire_con_out_stage6[187]), .inData_188(wire_con_out_stage6[188]), .inData_189(wire_con_out_stage6[189]), .inData_190(wire_con_out_stage6[190]), .inData_191(wire_con_out_stage6[191]), .inData_192(wire_con_out_stage6[192]), .inData_193(wire_con_out_stage6[193]), .inData_194(wire_con_out_stage6[194]), .inData_195(wire_con_out_stage6[195]), .inData_196(wire_con_out_stage6[196]), .inData_197(wire_con_out_stage6[197]), .inData_198(wire_con_out_stage6[198]), .inData_199(wire_con_out_stage6[199]), .inData_200(wire_con_out_stage6[200]), .inData_201(wire_con_out_stage6[201]), .inData_202(wire_con_out_stage6[202]), .inData_203(wire_con_out_stage6[203]), .inData_204(wire_con_out_stage6[204]), .inData_205(wire_con_out_stage6[205]), .inData_206(wire_con_out_stage6[206]), .inData_207(wire_con_out_stage6[207]), .inData_208(wire_con_out_stage6[208]), .inData_209(wire_con_out_stage6[209]), .inData_210(wire_con_out_stage6[210]), .inData_211(wire_con_out_stage6[211]), .inData_212(wire_con_out_stage6[212]), .inData_213(wire_con_out_stage6[213]), .inData_214(wire_con_out_stage6[214]), .inData_215(wire_con_out_stage6[215]), .inData_216(wire_con_out_stage6[216]), .inData_217(wire_con_out_stage6[217]), .inData_218(wire_con_out_stage6[218]), .inData_219(wire_con_out_stage6[219]), .inData_220(wire_con_out_stage6[220]), .inData_221(wire_con_out_stage6[221]), .inData_222(wire_con_out_stage6[222]), .inData_223(wire_con_out_stage6[223]), .inData_224(wire_con_out_stage6[224]), .inData_225(wire_con_out_stage6[225]), .inData_226(wire_con_out_stage6[226]), .inData_227(wire_con_out_stage6[227]), .inData_228(wire_con_out_stage6[228]), .inData_229(wire_con_out_stage6[229]), .inData_230(wire_con_out_stage6[230]), .inData_231(wire_con_out_stage6[231]), .inData_232(wire_con_out_stage6[232]), .inData_233(wire_con_out_stage6[233]), .inData_234(wire_con_out_stage6[234]), .inData_235(wire_con_out_stage6[235]), .inData_236(wire_con_out_stage6[236]), .inData_237(wire_con_out_stage6[237]), .inData_238(wire_con_out_stage6[238]), .inData_239(wire_con_out_stage6[239]), .inData_240(wire_con_out_stage6[240]), .inData_241(wire_con_out_stage6[241]), .inData_242(wire_con_out_stage6[242]), .inData_243(wire_con_out_stage6[243]), .inData_244(wire_con_out_stage6[244]), .inData_245(wire_con_out_stage6[245]), .inData_246(wire_con_out_stage6[246]), .inData_247(wire_con_out_stage6[247]), .inData_248(wire_con_out_stage6[248]), .inData_249(wire_con_out_stage6[249]), .inData_250(wire_con_out_stage6[250]), .inData_251(wire_con_out_stage6[251]), .inData_252(wire_con_out_stage6[252]), .inData_253(wire_con_out_stage6[253]), .inData_254(wire_con_out_stage6[254]), .inData_255(wire_con_out_stage6[255]), 
        .outData_0(wire_con_in_stage7[0]), .outData_1(wire_con_in_stage7[1]), .outData_2(wire_con_in_stage7[2]), .outData_3(wire_con_in_stage7[3]), .outData_4(wire_con_in_stage7[4]), .outData_5(wire_con_in_stage7[5]), .outData_6(wire_con_in_stage7[6]), .outData_7(wire_con_in_stage7[7]), .outData_8(wire_con_in_stage7[8]), .outData_9(wire_con_in_stage7[9]), .outData_10(wire_con_in_stage7[10]), .outData_11(wire_con_in_stage7[11]), .outData_12(wire_con_in_stage7[12]), .outData_13(wire_con_in_stage7[13]), .outData_14(wire_con_in_stage7[14]), .outData_15(wire_con_in_stage7[15]), .outData_16(wire_con_in_stage7[16]), .outData_17(wire_con_in_stage7[17]), .outData_18(wire_con_in_stage7[18]), .outData_19(wire_con_in_stage7[19]), .outData_20(wire_con_in_stage7[20]), .outData_21(wire_con_in_stage7[21]), .outData_22(wire_con_in_stage7[22]), .outData_23(wire_con_in_stage7[23]), .outData_24(wire_con_in_stage7[24]), .outData_25(wire_con_in_stage7[25]), .outData_26(wire_con_in_stage7[26]), .outData_27(wire_con_in_stage7[27]), .outData_28(wire_con_in_stage7[28]), .outData_29(wire_con_in_stage7[29]), .outData_30(wire_con_in_stage7[30]), .outData_31(wire_con_in_stage7[31]), .outData_32(wire_con_in_stage7[32]), .outData_33(wire_con_in_stage7[33]), .outData_34(wire_con_in_stage7[34]), .outData_35(wire_con_in_stage7[35]), .outData_36(wire_con_in_stage7[36]), .outData_37(wire_con_in_stage7[37]), .outData_38(wire_con_in_stage7[38]), .outData_39(wire_con_in_stage7[39]), .outData_40(wire_con_in_stage7[40]), .outData_41(wire_con_in_stage7[41]), .outData_42(wire_con_in_stage7[42]), .outData_43(wire_con_in_stage7[43]), .outData_44(wire_con_in_stage7[44]), .outData_45(wire_con_in_stage7[45]), .outData_46(wire_con_in_stage7[46]), .outData_47(wire_con_in_stage7[47]), .outData_48(wire_con_in_stage7[48]), .outData_49(wire_con_in_stage7[49]), .outData_50(wire_con_in_stage7[50]), .outData_51(wire_con_in_stage7[51]), .outData_52(wire_con_in_stage7[52]), .outData_53(wire_con_in_stage7[53]), .outData_54(wire_con_in_stage7[54]), .outData_55(wire_con_in_stage7[55]), .outData_56(wire_con_in_stage7[56]), .outData_57(wire_con_in_stage7[57]), .outData_58(wire_con_in_stage7[58]), .outData_59(wire_con_in_stage7[59]), .outData_60(wire_con_in_stage7[60]), .outData_61(wire_con_in_stage7[61]), .outData_62(wire_con_in_stage7[62]), .outData_63(wire_con_in_stage7[63]), .outData_64(wire_con_in_stage7[64]), .outData_65(wire_con_in_stage7[65]), .outData_66(wire_con_in_stage7[66]), .outData_67(wire_con_in_stage7[67]), .outData_68(wire_con_in_stage7[68]), .outData_69(wire_con_in_stage7[69]), .outData_70(wire_con_in_stage7[70]), .outData_71(wire_con_in_stage7[71]), .outData_72(wire_con_in_stage7[72]), .outData_73(wire_con_in_stage7[73]), .outData_74(wire_con_in_stage7[74]), .outData_75(wire_con_in_stage7[75]), .outData_76(wire_con_in_stage7[76]), .outData_77(wire_con_in_stage7[77]), .outData_78(wire_con_in_stage7[78]), .outData_79(wire_con_in_stage7[79]), .outData_80(wire_con_in_stage7[80]), .outData_81(wire_con_in_stage7[81]), .outData_82(wire_con_in_stage7[82]), .outData_83(wire_con_in_stage7[83]), .outData_84(wire_con_in_stage7[84]), .outData_85(wire_con_in_stage7[85]), .outData_86(wire_con_in_stage7[86]), .outData_87(wire_con_in_stage7[87]), .outData_88(wire_con_in_stage7[88]), .outData_89(wire_con_in_stage7[89]), .outData_90(wire_con_in_stage7[90]), .outData_91(wire_con_in_stage7[91]), .outData_92(wire_con_in_stage7[92]), .outData_93(wire_con_in_stage7[93]), .outData_94(wire_con_in_stage7[94]), .outData_95(wire_con_in_stage7[95]), .outData_96(wire_con_in_stage7[96]), .outData_97(wire_con_in_stage7[97]), .outData_98(wire_con_in_stage7[98]), .outData_99(wire_con_in_stage7[99]), .outData_100(wire_con_in_stage7[100]), .outData_101(wire_con_in_stage7[101]), .outData_102(wire_con_in_stage7[102]), .outData_103(wire_con_in_stage7[103]), .outData_104(wire_con_in_stage7[104]), .outData_105(wire_con_in_stage7[105]), .outData_106(wire_con_in_stage7[106]), .outData_107(wire_con_in_stage7[107]), .outData_108(wire_con_in_stage7[108]), .outData_109(wire_con_in_stage7[109]), .outData_110(wire_con_in_stage7[110]), .outData_111(wire_con_in_stage7[111]), .outData_112(wire_con_in_stage7[112]), .outData_113(wire_con_in_stage7[113]), .outData_114(wire_con_in_stage7[114]), .outData_115(wire_con_in_stage7[115]), .outData_116(wire_con_in_stage7[116]), .outData_117(wire_con_in_stage7[117]), .outData_118(wire_con_in_stage7[118]), .outData_119(wire_con_in_stage7[119]), .outData_120(wire_con_in_stage7[120]), .outData_121(wire_con_in_stage7[121]), .outData_122(wire_con_in_stage7[122]), .outData_123(wire_con_in_stage7[123]), .outData_124(wire_con_in_stage7[124]), .outData_125(wire_con_in_stage7[125]), .outData_126(wire_con_in_stage7[126]), .outData_127(wire_con_in_stage7[127]), .outData_128(wire_con_in_stage7[128]), .outData_129(wire_con_in_stage7[129]), .outData_130(wire_con_in_stage7[130]), .outData_131(wire_con_in_stage7[131]), .outData_132(wire_con_in_stage7[132]), .outData_133(wire_con_in_stage7[133]), .outData_134(wire_con_in_stage7[134]), .outData_135(wire_con_in_stage7[135]), .outData_136(wire_con_in_stage7[136]), .outData_137(wire_con_in_stage7[137]), .outData_138(wire_con_in_stage7[138]), .outData_139(wire_con_in_stage7[139]), .outData_140(wire_con_in_stage7[140]), .outData_141(wire_con_in_stage7[141]), .outData_142(wire_con_in_stage7[142]), .outData_143(wire_con_in_stage7[143]), .outData_144(wire_con_in_stage7[144]), .outData_145(wire_con_in_stage7[145]), .outData_146(wire_con_in_stage7[146]), .outData_147(wire_con_in_stage7[147]), .outData_148(wire_con_in_stage7[148]), .outData_149(wire_con_in_stage7[149]), .outData_150(wire_con_in_stage7[150]), .outData_151(wire_con_in_stage7[151]), .outData_152(wire_con_in_stage7[152]), .outData_153(wire_con_in_stage7[153]), .outData_154(wire_con_in_stage7[154]), .outData_155(wire_con_in_stage7[155]), .outData_156(wire_con_in_stage7[156]), .outData_157(wire_con_in_stage7[157]), .outData_158(wire_con_in_stage7[158]), .outData_159(wire_con_in_stage7[159]), .outData_160(wire_con_in_stage7[160]), .outData_161(wire_con_in_stage7[161]), .outData_162(wire_con_in_stage7[162]), .outData_163(wire_con_in_stage7[163]), .outData_164(wire_con_in_stage7[164]), .outData_165(wire_con_in_stage7[165]), .outData_166(wire_con_in_stage7[166]), .outData_167(wire_con_in_stage7[167]), .outData_168(wire_con_in_stage7[168]), .outData_169(wire_con_in_stage7[169]), .outData_170(wire_con_in_stage7[170]), .outData_171(wire_con_in_stage7[171]), .outData_172(wire_con_in_stage7[172]), .outData_173(wire_con_in_stage7[173]), .outData_174(wire_con_in_stage7[174]), .outData_175(wire_con_in_stage7[175]), .outData_176(wire_con_in_stage7[176]), .outData_177(wire_con_in_stage7[177]), .outData_178(wire_con_in_stage7[178]), .outData_179(wire_con_in_stage7[179]), .outData_180(wire_con_in_stage7[180]), .outData_181(wire_con_in_stage7[181]), .outData_182(wire_con_in_stage7[182]), .outData_183(wire_con_in_stage7[183]), .outData_184(wire_con_in_stage7[184]), .outData_185(wire_con_in_stage7[185]), .outData_186(wire_con_in_stage7[186]), .outData_187(wire_con_in_stage7[187]), .outData_188(wire_con_in_stage7[188]), .outData_189(wire_con_in_stage7[189]), .outData_190(wire_con_in_stage7[190]), .outData_191(wire_con_in_stage7[191]), .outData_192(wire_con_in_stage7[192]), .outData_193(wire_con_in_stage7[193]), .outData_194(wire_con_in_stage7[194]), .outData_195(wire_con_in_stage7[195]), .outData_196(wire_con_in_stage7[196]), .outData_197(wire_con_in_stage7[197]), .outData_198(wire_con_in_stage7[198]), .outData_199(wire_con_in_stage7[199]), .outData_200(wire_con_in_stage7[200]), .outData_201(wire_con_in_stage7[201]), .outData_202(wire_con_in_stage7[202]), .outData_203(wire_con_in_stage7[203]), .outData_204(wire_con_in_stage7[204]), .outData_205(wire_con_in_stage7[205]), .outData_206(wire_con_in_stage7[206]), .outData_207(wire_con_in_stage7[207]), .outData_208(wire_con_in_stage7[208]), .outData_209(wire_con_in_stage7[209]), .outData_210(wire_con_in_stage7[210]), .outData_211(wire_con_in_stage7[211]), .outData_212(wire_con_in_stage7[212]), .outData_213(wire_con_in_stage7[213]), .outData_214(wire_con_in_stage7[214]), .outData_215(wire_con_in_stage7[215]), .outData_216(wire_con_in_stage7[216]), .outData_217(wire_con_in_stage7[217]), .outData_218(wire_con_in_stage7[218]), .outData_219(wire_con_in_stage7[219]), .outData_220(wire_con_in_stage7[220]), .outData_221(wire_con_in_stage7[221]), .outData_222(wire_con_in_stage7[222]), .outData_223(wire_con_in_stage7[223]), .outData_224(wire_con_in_stage7[224]), .outData_225(wire_con_in_stage7[225]), .outData_226(wire_con_in_stage7[226]), .outData_227(wire_con_in_stage7[227]), .outData_228(wire_con_in_stage7[228]), .outData_229(wire_con_in_stage7[229]), .outData_230(wire_con_in_stage7[230]), .outData_231(wire_con_in_stage7[231]), .outData_232(wire_con_in_stage7[232]), .outData_233(wire_con_in_stage7[233]), .outData_234(wire_con_in_stage7[234]), .outData_235(wire_con_in_stage7[235]), .outData_236(wire_con_in_stage7[236]), .outData_237(wire_con_in_stage7[237]), .outData_238(wire_con_in_stage7[238]), .outData_239(wire_con_in_stage7[239]), .outData_240(wire_con_in_stage7[240]), .outData_241(wire_con_in_stage7[241]), .outData_242(wire_con_in_stage7[242]), .outData_243(wire_con_in_stage7[243]), .outData_244(wire_con_in_stage7[244]), .outData_245(wire_con_in_stage7[245]), .outData_246(wire_con_in_stage7[246]), .outData_247(wire_con_in_stage7[247]), .outData_248(wire_con_in_stage7[248]), .outData_249(wire_con_in_stage7[249]), .outData_250(wire_con_in_stage7[250]), .outData_251(wire_con_in_stage7[251]), .outData_252(wire_con_in_stage7[252]), .outData_253(wire_con_in_stage7[253]), .outData_254(wire_con_in_stage7[254]), .outData_255(wire_con_in_stage7[255]), 
        .in_start(in_start_stage7), .out_start(con_in_start_stage7), .ctrl(wire_ctrl_stage7), .clk(clk), .rst(rst));
  
  wireCon_dp256_st7_L wire_stage_7(
        .inData_0(wire_con_in_stage7[0]), .inData_1(wire_con_in_stage7[1]), .inData_2(wire_con_in_stage7[2]), .inData_3(wire_con_in_stage7[3]), .inData_4(wire_con_in_stage7[4]), .inData_5(wire_con_in_stage7[5]), .inData_6(wire_con_in_stage7[6]), .inData_7(wire_con_in_stage7[7]), .inData_8(wire_con_in_stage7[8]), .inData_9(wire_con_in_stage7[9]), .inData_10(wire_con_in_stage7[10]), .inData_11(wire_con_in_stage7[11]), .inData_12(wire_con_in_stage7[12]), .inData_13(wire_con_in_stage7[13]), .inData_14(wire_con_in_stage7[14]), .inData_15(wire_con_in_stage7[15]), .inData_16(wire_con_in_stage7[16]), .inData_17(wire_con_in_stage7[17]), .inData_18(wire_con_in_stage7[18]), .inData_19(wire_con_in_stage7[19]), .inData_20(wire_con_in_stage7[20]), .inData_21(wire_con_in_stage7[21]), .inData_22(wire_con_in_stage7[22]), .inData_23(wire_con_in_stage7[23]), .inData_24(wire_con_in_stage7[24]), .inData_25(wire_con_in_stage7[25]), .inData_26(wire_con_in_stage7[26]), .inData_27(wire_con_in_stage7[27]), .inData_28(wire_con_in_stage7[28]), .inData_29(wire_con_in_stage7[29]), .inData_30(wire_con_in_stage7[30]), .inData_31(wire_con_in_stage7[31]), .inData_32(wire_con_in_stage7[32]), .inData_33(wire_con_in_stage7[33]), .inData_34(wire_con_in_stage7[34]), .inData_35(wire_con_in_stage7[35]), .inData_36(wire_con_in_stage7[36]), .inData_37(wire_con_in_stage7[37]), .inData_38(wire_con_in_stage7[38]), .inData_39(wire_con_in_stage7[39]), .inData_40(wire_con_in_stage7[40]), .inData_41(wire_con_in_stage7[41]), .inData_42(wire_con_in_stage7[42]), .inData_43(wire_con_in_stage7[43]), .inData_44(wire_con_in_stage7[44]), .inData_45(wire_con_in_stage7[45]), .inData_46(wire_con_in_stage7[46]), .inData_47(wire_con_in_stage7[47]), .inData_48(wire_con_in_stage7[48]), .inData_49(wire_con_in_stage7[49]), .inData_50(wire_con_in_stage7[50]), .inData_51(wire_con_in_stage7[51]), .inData_52(wire_con_in_stage7[52]), .inData_53(wire_con_in_stage7[53]), .inData_54(wire_con_in_stage7[54]), .inData_55(wire_con_in_stage7[55]), .inData_56(wire_con_in_stage7[56]), .inData_57(wire_con_in_stage7[57]), .inData_58(wire_con_in_stage7[58]), .inData_59(wire_con_in_stage7[59]), .inData_60(wire_con_in_stage7[60]), .inData_61(wire_con_in_stage7[61]), .inData_62(wire_con_in_stage7[62]), .inData_63(wire_con_in_stage7[63]), .inData_64(wire_con_in_stage7[64]), .inData_65(wire_con_in_stage7[65]), .inData_66(wire_con_in_stage7[66]), .inData_67(wire_con_in_stage7[67]), .inData_68(wire_con_in_stage7[68]), .inData_69(wire_con_in_stage7[69]), .inData_70(wire_con_in_stage7[70]), .inData_71(wire_con_in_stage7[71]), .inData_72(wire_con_in_stage7[72]), .inData_73(wire_con_in_stage7[73]), .inData_74(wire_con_in_stage7[74]), .inData_75(wire_con_in_stage7[75]), .inData_76(wire_con_in_stage7[76]), .inData_77(wire_con_in_stage7[77]), .inData_78(wire_con_in_stage7[78]), .inData_79(wire_con_in_stage7[79]), .inData_80(wire_con_in_stage7[80]), .inData_81(wire_con_in_stage7[81]), .inData_82(wire_con_in_stage7[82]), .inData_83(wire_con_in_stage7[83]), .inData_84(wire_con_in_stage7[84]), .inData_85(wire_con_in_stage7[85]), .inData_86(wire_con_in_stage7[86]), .inData_87(wire_con_in_stage7[87]), .inData_88(wire_con_in_stage7[88]), .inData_89(wire_con_in_stage7[89]), .inData_90(wire_con_in_stage7[90]), .inData_91(wire_con_in_stage7[91]), .inData_92(wire_con_in_stage7[92]), .inData_93(wire_con_in_stage7[93]), .inData_94(wire_con_in_stage7[94]), .inData_95(wire_con_in_stage7[95]), .inData_96(wire_con_in_stage7[96]), .inData_97(wire_con_in_stage7[97]), .inData_98(wire_con_in_stage7[98]), .inData_99(wire_con_in_stage7[99]), .inData_100(wire_con_in_stage7[100]), .inData_101(wire_con_in_stage7[101]), .inData_102(wire_con_in_stage7[102]), .inData_103(wire_con_in_stage7[103]), .inData_104(wire_con_in_stage7[104]), .inData_105(wire_con_in_stage7[105]), .inData_106(wire_con_in_stage7[106]), .inData_107(wire_con_in_stage7[107]), .inData_108(wire_con_in_stage7[108]), .inData_109(wire_con_in_stage7[109]), .inData_110(wire_con_in_stage7[110]), .inData_111(wire_con_in_stage7[111]), .inData_112(wire_con_in_stage7[112]), .inData_113(wire_con_in_stage7[113]), .inData_114(wire_con_in_stage7[114]), .inData_115(wire_con_in_stage7[115]), .inData_116(wire_con_in_stage7[116]), .inData_117(wire_con_in_stage7[117]), .inData_118(wire_con_in_stage7[118]), .inData_119(wire_con_in_stage7[119]), .inData_120(wire_con_in_stage7[120]), .inData_121(wire_con_in_stage7[121]), .inData_122(wire_con_in_stage7[122]), .inData_123(wire_con_in_stage7[123]), .inData_124(wire_con_in_stage7[124]), .inData_125(wire_con_in_stage7[125]), .inData_126(wire_con_in_stage7[126]), .inData_127(wire_con_in_stage7[127]), .inData_128(wire_con_in_stage7[128]), .inData_129(wire_con_in_stage7[129]), .inData_130(wire_con_in_stage7[130]), .inData_131(wire_con_in_stage7[131]), .inData_132(wire_con_in_stage7[132]), .inData_133(wire_con_in_stage7[133]), .inData_134(wire_con_in_stage7[134]), .inData_135(wire_con_in_stage7[135]), .inData_136(wire_con_in_stage7[136]), .inData_137(wire_con_in_stage7[137]), .inData_138(wire_con_in_stage7[138]), .inData_139(wire_con_in_stage7[139]), .inData_140(wire_con_in_stage7[140]), .inData_141(wire_con_in_stage7[141]), .inData_142(wire_con_in_stage7[142]), .inData_143(wire_con_in_stage7[143]), .inData_144(wire_con_in_stage7[144]), .inData_145(wire_con_in_stage7[145]), .inData_146(wire_con_in_stage7[146]), .inData_147(wire_con_in_stage7[147]), .inData_148(wire_con_in_stage7[148]), .inData_149(wire_con_in_stage7[149]), .inData_150(wire_con_in_stage7[150]), .inData_151(wire_con_in_stage7[151]), .inData_152(wire_con_in_stage7[152]), .inData_153(wire_con_in_stage7[153]), .inData_154(wire_con_in_stage7[154]), .inData_155(wire_con_in_stage7[155]), .inData_156(wire_con_in_stage7[156]), .inData_157(wire_con_in_stage7[157]), .inData_158(wire_con_in_stage7[158]), .inData_159(wire_con_in_stage7[159]), .inData_160(wire_con_in_stage7[160]), .inData_161(wire_con_in_stage7[161]), .inData_162(wire_con_in_stage7[162]), .inData_163(wire_con_in_stage7[163]), .inData_164(wire_con_in_stage7[164]), .inData_165(wire_con_in_stage7[165]), .inData_166(wire_con_in_stage7[166]), .inData_167(wire_con_in_stage7[167]), .inData_168(wire_con_in_stage7[168]), .inData_169(wire_con_in_stage7[169]), .inData_170(wire_con_in_stage7[170]), .inData_171(wire_con_in_stage7[171]), .inData_172(wire_con_in_stage7[172]), .inData_173(wire_con_in_stage7[173]), .inData_174(wire_con_in_stage7[174]), .inData_175(wire_con_in_stage7[175]), .inData_176(wire_con_in_stage7[176]), .inData_177(wire_con_in_stage7[177]), .inData_178(wire_con_in_stage7[178]), .inData_179(wire_con_in_stage7[179]), .inData_180(wire_con_in_stage7[180]), .inData_181(wire_con_in_stage7[181]), .inData_182(wire_con_in_stage7[182]), .inData_183(wire_con_in_stage7[183]), .inData_184(wire_con_in_stage7[184]), .inData_185(wire_con_in_stage7[185]), .inData_186(wire_con_in_stage7[186]), .inData_187(wire_con_in_stage7[187]), .inData_188(wire_con_in_stage7[188]), .inData_189(wire_con_in_stage7[189]), .inData_190(wire_con_in_stage7[190]), .inData_191(wire_con_in_stage7[191]), .inData_192(wire_con_in_stage7[192]), .inData_193(wire_con_in_stage7[193]), .inData_194(wire_con_in_stage7[194]), .inData_195(wire_con_in_stage7[195]), .inData_196(wire_con_in_stage7[196]), .inData_197(wire_con_in_stage7[197]), .inData_198(wire_con_in_stage7[198]), .inData_199(wire_con_in_stage7[199]), .inData_200(wire_con_in_stage7[200]), .inData_201(wire_con_in_stage7[201]), .inData_202(wire_con_in_stage7[202]), .inData_203(wire_con_in_stage7[203]), .inData_204(wire_con_in_stage7[204]), .inData_205(wire_con_in_stage7[205]), .inData_206(wire_con_in_stage7[206]), .inData_207(wire_con_in_stage7[207]), .inData_208(wire_con_in_stage7[208]), .inData_209(wire_con_in_stage7[209]), .inData_210(wire_con_in_stage7[210]), .inData_211(wire_con_in_stage7[211]), .inData_212(wire_con_in_stage7[212]), .inData_213(wire_con_in_stage7[213]), .inData_214(wire_con_in_stage7[214]), .inData_215(wire_con_in_stage7[215]), .inData_216(wire_con_in_stage7[216]), .inData_217(wire_con_in_stage7[217]), .inData_218(wire_con_in_stage7[218]), .inData_219(wire_con_in_stage7[219]), .inData_220(wire_con_in_stage7[220]), .inData_221(wire_con_in_stage7[221]), .inData_222(wire_con_in_stage7[222]), .inData_223(wire_con_in_stage7[223]), .inData_224(wire_con_in_stage7[224]), .inData_225(wire_con_in_stage7[225]), .inData_226(wire_con_in_stage7[226]), .inData_227(wire_con_in_stage7[227]), .inData_228(wire_con_in_stage7[228]), .inData_229(wire_con_in_stage7[229]), .inData_230(wire_con_in_stage7[230]), .inData_231(wire_con_in_stage7[231]), .inData_232(wire_con_in_stage7[232]), .inData_233(wire_con_in_stage7[233]), .inData_234(wire_con_in_stage7[234]), .inData_235(wire_con_in_stage7[235]), .inData_236(wire_con_in_stage7[236]), .inData_237(wire_con_in_stage7[237]), .inData_238(wire_con_in_stage7[238]), .inData_239(wire_con_in_stage7[239]), .inData_240(wire_con_in_stage7[240]), .inData_241(wire_con_in_stage7[241]), .inData_242(wire_con_in_stage7[242]), .inData_243(wire_con_in_stage7[243]), .inData_244(wire_con_in_stage7[244]), .inData_245(wire_con_in_stage7[245]), .inData_246(wire_con_in_stage7[246]), .inData_247(wire_con_in_stage7[247]), .inData_248(wire_con_in_stage7[248]), .inData_249(wire_con_in_stage7[249]), .inData_250(wire_con_in_stage7[250]), .inData_251(wire_con_in_stage7[251]), .inData_252(wire_con_in_stage7[252]), .inData_253(wire_con_in_stage7[253]), .inData_254(wire_con_in_stage7[254]), .inData_255(wire_con_in_stage7[255]), 
        .outData_0(wireOut[0]), .outData_1(wireOut[1]), .outData_2(wireOut[2]), .outData_3(wireOut[3]), .outData_4(wireOut[4]), .outData_5(wireOut[5]), .outData_6(wireOut[6]), .outData_7(wireOut[7]), .outData_8(wireOut[8]), .outData_9(wireOut[9]), .outData_10(wireOut[10]), .outData_11(wireOut[11]), .outData_12(wireOut[12]), .outData_13(wireOut[13]), .outData_14(wireOut[14]), .outData_15(wireOut[15]), .outData_16(wireOut[16]), .outData_17(wireOut[17]), .outData_18(wireOut[18]), .outData_19(wireOut[19]), .outData_20(wireOut[20]), .outData_21(wireOut[21]), .outData_22(wireOut[22]), .outData_23(wireOut[23]), .outData_24(wireOut[24]), .outData_25(wireOut[25]), .outData_26(wireOut[26]), .outData_27(wireOut[27]), .outData_28(wireOut[28]), .outData_29(wireOut[29]), .outData_30(wireOut[30]), .outData_31(wireOut[31]), .outData_32(wireOut[32]), .outData_33(wireOut[33]), .outData_34(wireOut[34]), .outData_35(wireOut[35]), .outData_36(wireOut[36]), .outData_37(wireOut[37]), .outData_38(wireOut[38]), .outData_39(wireOut[39]), .outData_40(wireOut[40]), .outData_41(wireOut[41]), .outData_42(wireOut[42]), .outData_43(wireOut[43]), .outData_44(wireOut[44]), .outData_45(wireOut[45]), .outData_46(wireOut[46]), .outData_47(wireOut[47]), .outData_48(wireOut[48]), .outData_49(wireOut[49]), .outData_50(wireOut[50]), .outData_51(wireOut[51]), .outData_52(wireOut[52]), .outData_53(wireOut[53]), .outData_54(wireOut[54]), .outData_55(wireOut[55]), .outData_56(wireOut[56]), .outData_57(wireOut[57]), .outData_58(wireOut[58]), .outData_59(wireOut[59]), .outData_60(wireOut[60]), .outData_61(wireOut[61]), .outData_62(wireOut[62]), .outData_63(wireOut[63]), .outData_64(wireOut[64]), .outData_65(wireOut[65]), .outData_66(wireOut[66]), .outData_67(wireOut[67]), .outData_68(wireOut[68]), .outData_69(wireOut[69]), .outData_70(wireOut[70]), .outData_71(wireOut[71]), .outData_72(wireOut[72]), .outData_73(wireOut[73]), .outData_74(wireOut[74]), .outData_75(wireOut[75]), .outData_76(wireOut[76]), .outData_77(wireOut[77]), .outData_78(wireOut[78]), .outData_79(wireOut[79]), .outData_80(wireOut[80]), .outData_81(wireOut[81]), .outData_82(wireOut[82]), .outData_83(wireOut[83]), .outData_84(wireOut[84]), .outData_85(wireOut[85]), .outData_86(wireOut[86]), .outData_87(wireOut[87]), .outData_88(wireOut[88]), .outData_89(wireOut[89]), .outData_90(wireOut[90]), .outData_91(wireOut[91]), .outData_92(wireOut[92]), .outData_93(wireOut[93]), .outData_94(wireOut[94]), .outData_95(wireOut[95]), .outData_96(wireOut[96]), .outData_97(wireOut[97]), .outData_98(wireOut[98]), .outData_99(wireOut[99]), .outData_100(wireOut[100]), .outData_101(wireOut[101]), .outData_102(wireOut[102]), .outData_103(wireOut[103]), .outData_104(wireOut[104]), .outData_105(wireOut[105]), .outData_106(wireOut[106]), .outData_107(wireOut[107]), .outData_108(wireOut[108]), .outData_109(wireOut[109]), .outData_110(wireOut[110]), .outData_111(wireOut[111]), .outData_112(wireOut[112]), .outData_113(wireOut[113]), .outData_114(wireOut[114]), .outData_115(wireOut[115]), .outData_116(wireOut[116]), .outData_117(wireOut[117]), .outData_118(wireOut[118]), .outData_119(wireOut[119]), .outData_120(wireOut[120]), .outData_121(wireOut[121]), .outData_122(wireOut[122]), .outData_123(wireOut[123]), .outData_124(wireOut[124]), .outData_125(wireOut[125]), .outData_126(wireOut[126]), .outData_127(wireOut[127]), .outData_128(wireOut[128]), .outData_129(wireOut[129]), .outData_130(wireOut[130]), .outData_131(wireOut[131]), .outData_132(wireOut[132]), .outData_133(wireOut[133]), .outData_134(wireOut[134]), .outData_135(wireOut[135]), .outData_136(wireOut[136]), .outData_137(wireOut[137]), .outData_138(wireOut[138]), .outData_139(wireOut[139]), .outData_140(wireOut[140]), .outData_141(wireOut[141]), .outData_142(wireOut[142]), .outData_143(wireOut[143]), .outData_144(wireOut[144]), .outData_145(wireOut[145]), .outData_146(wireOut[146]), .outData_147(wireOut[147]), .outData_148(wireOut[148]), .outData_149(wireOut[149]), .outData_150(wireOut[150]), .outData_151(wireOut[151]), .outData_152(wireOut[152]), .outData_153(wireOut[153]), .outData_154(wireOut[154]), .outData_155(wireOut[155]), .outData_156(wireOut[156]), .outData_157(wireOut[157]), .outData_158(wireOut[158]), .outData_159(wireOut[159]), .outData_160(wireOut[160]), .outData_161(wireOut[161]), .outData_162(wireOut[162]), .outData_163(wireOut[163]), .outData_164(wireOut[164]), .outData_165(wireOut[165]), .outData_166(wireOut[166]), .outData_167(wireOut[167]), .outData_168(wireOut[168]), .outData_169(wireOut[169]), .outData_170(wireOut[170]), .outData_171(wireOut[171]), .outData_172(wireOut[172]), .outData_173(wireOut[173]), .outData_174(wireOut[174]), .outData_175(wireOut[175]), .outData_176(wireOut[176]), .outData_177(wireOut[177]), .outData_178(wireOut[178]), .outData_179(wireOut[179]), .outData_180(wireOut[180]), .outData_181(wireOut[181]), .outData_182(wireOut[182]), .outData_183(wireOut[183]), .outData_184(wireOut[184]), .outData_185(wireOut[185]), .outData_186(wireOut[186]), .outData_187(wireOut[187]), .outData_188(wireOut[188]), .outData_189(wireOut[189]), .outData_190(wireOut[190]), .outData_191(wireOut[191]), .outData_192(wireOut[192]), .outData_193(wireOut[193]), .outData_194(wireOut[194]), .outData_195(wireOut[195]), .outData_196(wireOut[196]), .outData_197(wireOut[197]), .outData_198(wireOut[198]), .outData_199(wireOut[199]), .outData_200(wireOut[200]), .outData_201(wireOut[201]), .outData_202(wireOut[202]), .outData_203(wireOut[203]), .outData_204(wireOut[204]), .outData_205(wireOut[205]), .outData_206(wireOut[206]), .outData_207(wireOut[207]), .outData_208(wireOut[208]), .outData_209(wireOut[209]), .outData_210(wireOut[210]), .outData_211(wireOut[211]), .outData_212(wireOut[212]), .outData_213(wireOut[213]), .outData_214(wireOut[214]), .outData_215(wireOut[215]), .outData_216(wireOut[216]), .outData_217(wireOut[217]), .outData_218(wireOut[218]), .outData_219(wireOut[219]), .outData_220(wireOut[220]), .outData_221(wireOut[221]), .outData_222(wireOut[222]), .outData_223(wireOut[223]), .outData_224(wireOut[224]), .outData_225(wireOut[225]), .outData_226(wireOut[226]), .outData_227(wireOut[227]), .outData_228(wireOut[228]), .outData_229(wireOut[229]), .outData_230(wireOut[230]), .outData_231(wireOut[231]), .outData_232(wireOut[232]), .outData_233(wireOut[233]), .outData_234(wireOut[234]), .outData_235(wireOut[235]), .outData_236(wireOut[236]), .outData_237(wireOut[237]), .outData_238(wireOut[238]), .outData_239(wireOut[239]), .outData_240(wireOut[240]), .outData_241(wireOut[241]), .outData_242(wireOut[242]), .outData_243(wireOut[243]), .outData_244(wireOut[244]), .outData_245(wireOut[245]), .outData_246(wireOut[246]), .outData_247(wireOut[247]), .outData_248(wireOut[248]), .outData_249(wireOut[249]), .outData_250(wireOut[250]), .outData_251(wireOut[251]), .outData_252(wireOut[252]), .outData_253(wireOut[253]), .outData_254(wireOut[254]), .outData_255(wireOut[255]), 
        .in_start(con_in_start_stage7), .out_start(out_start_w), .clk(clk), .rst(rst)); 

  
  assign wire_ctrl_stage7[0] = counter_w[0]; 
  assign wire_ctrl_stage7[1] = counter_w[0]; 
  assign wire_ctrl_stage7[2] = counter_w[0]; 
  assign wire_ctrl_stage7[3] = counter_w[0]; 
  assign wire_ctrl_stage7[4] = counter_w[0]; 
  assign wire_ctrl_stage7[5] = counter_w[0]; 
  assign wire_ctrl_stage7[6] = counter_w[0]; 
  assign wire_ctrl_stage7[7] = counter_w[0]; 
  assign wire_ctrl_stage7[8] = counter_w[0]; 
  assign wire_ctrl_stage7[9] = counter_w[0]; 
  assign wire_ctrl_stage7[10] = counter_w[0]; 
  assign wire_ctrl_stage7[11] = counter_w[0]; 
  assign wire_ctrl_stage7[12] = counter_w[0]; 
  assign wire_ctrl_stage7[13] = counter_w[0]; 
  assign wire_ctrl_stage7[14] = counter_w[0]; 
  assign wire_ctrl_stage7[15] = counter_w[0]; 
  assign wire_ctrl_stage7[16] = counter_w[0]; 
  assign wire_ctrl_stage7[17] = counter_w[0]; 
  assign wire_ctrl_stage7[18] = counter_w[0]; 
  assign wire_ctrl_stage7[19] = counter_w[0]; 
  assign wire_ctrl_stage7[20] = counter_w[0]; 
  assign wire_ctrl_stage7[21] = counter_w[0]; 
  assign wire_ctrl_stage7[22] = counter_w[0]; 
  assign wire_ctrl_stage7[23] = counter_w[0]; 
  assign wire_ctrl_stage7[24] = counter_w[0]; 
  assign wire_ctrl_stage7[25] = counter_w[0]; 
  assign wire_ctrl_stage7[26] = counter_w[0]; 
  assign wire_ctrl_stage7[27] = counter_w[0]; 
  assign wire_ctrl_stage7[28] = counter_w[0]; 
  assign wire_ctrl_stage7[29] = counter_w[0]; 
  assign wire_ctrl_stage7[30] = counter_w[0]; 
  assign wire_ctrl_stage7[31] = counter_w[0]; 
  assign wire_ctrl_stage7[32] = counter_w[0]; 
  assign wire_ctrl_stage7[33] = counter_w[0]; 
  assign wire_ctrl_stage7[34] = counter_w[0]; 
  assign wire_ctrl_stage7[35] = counter_w[0]; 
  assign wire_ctrl_stage7[36] = counter_w[0]; 
  assign wire_ctrl_stage7[37] = counter_w[0]; 
  assign wire_ctrl_stage7[38] = counter_w[0]; 
  assign wire_ctrl_stage7[39] = counter_w[0]; 
  assign wire_ctrl_stage7[40] = counter_w[0]; 
  assign wire_ctrl_stage7[41] = counter_w[0]; 
  assign wire_ctrl_stage7[42] = counter_w[0]; 
  assign wire_ctrl_stage7[43] = counter_w[0]; 
  assign wire_ctrl_stage7[44] = counter_w[0]; 
  assign wire_ctrl_stage7[45] = counter_w[0]; 
  assign wire_ctrl_stage7[46] = counter_w[0]; 
  assign wire_ctrl_stage7[47] = counter_w[0]; 
  assign wire_ctrl_stage7[48] = counter_w[0]; 
  assign wire_ctrl_stage7[49] = counter_w[0]; 
  assign wire_ctrl_stage7[50] = counter_w[0]; 
  assign wire_ctrl_stage7[51] = counter_w[0]; 
  assign wire_ctrl_stage7[52] = counter_w[0]; 
  assign wire_ctrl_stage7[53] = counter_w[0]; 
  assign wire_ctrl_stage7[54] = counter_w[0]; 
  assign wire_ctrl_stage7[55] = counter_w[0]; 
  assign wire_ctrl_stage7[56] = counter_w[0]; 
  assign wire_ctrl_stage7[57] = counter_w[0]; 
  assign wire_ctrl_stage7[58] = counter_w[0]; 
  assign wire_ctrl_stage7[59] = counter_w[0]; 
  assign wire_ctrl_stage7[60] = counter_w[0]; 
  assign wire_ctrl_stage7[61] = counter_w[0]; 
  assign wire_ctrl_stage7[62] = counter_w[0]; 
  assign wire_ctrl_stage7[63] = counter_w[0]; 
  assign wire_ctrl_stage7[64] = counter_w[0]; 
  assign wire_ctrl_stage7[65] = counter_w[0]; 
  assign wire_ctrl_stage7[66] = counter_w[0]; 
  assign wire_ctrl_stage7[67] = counter_w[0]; 
  assign wire_ctrl_stage7[68] = counter_w[0]; 
  assign wire_ctrl_stage7[69] = counter_w[0]; 
  assign wire_ctrl_stage7[70] = counter_w[0]; 
  assign wire_ctrl_stage7[71] = counter_w[0]; 
  assign wire_ctrl_stage7[72] = counter_w[0]; 
  assign wire_ctrl_stage7[73] = counter_w[0]; 
  assign wire_ctrl_stage7[74] = counter_w[0]; 
  assign wire_ctrl_stage7[75] = counter_w[0]; 
  assign wire_ctrl_stage7[76] = counter_w[0]; 
  assign wire_ctrl_stage7[77] = counter_w[0]; 
  assign wire_ctrl_stage7[78] = counter_w[0]; 
  assign wire_ctrl_stage7[79] = counter_w[0]; 
  assign wire_ctrl_stage7[80] = counter_w[0]; 
  assign wire_ctrl_stage7[81] = counter_w[0]; 
  assign wire_ctrl_stage7[82] = counter_w[0]; 
  assign wire_ctrl_stage7[83] = counter_w[0]; 
  assign wire_ctrl_stage7[84] = counter_w[0]; 
  assign wire_ctrl_stage7[85] = counter_w[0]; 
  assign wire_ctrl_stage7[86] = counter_w[0]; 
  assign wire_ctrl_stage7[87] = counter_w[0]; 
  assign wire_ctrl_stage7[88] = counter_w[0]; 
  assign wire_ctrl_stage7[89] = counter_w[0]; 
  assign wire_ctrl_stage7[90] = counter_w[0]; 
  assign wire_ctrl_stage7[91] = counter_w[0]; 
  assign wire_ctrl_stage7[92] = counter_w[0]; 
  assign wire_ctrl_stage7[93] = counter_w[0]; 
  assign wire_ctrl_stage7[94] = counter_w[0]; 
  assign wire_ctrl_stage7[95] = counter_w[0]; 
  assign wire_ctrl_stage7[96] = counter_w[0]; 
  assign wire_ctrl_stage7[97] = counter_w[0]; 
  assign wire_ctrl_stage7[98] = counter_w[0]; 
  assign wire_ctrl_stage7[99] = counter_w[0]; 
  assign wire_ctrl_stage7[100] = counter_w[0]; 
  assign wire_ctrl_stage7[101] = counter_w[0]; 
  assign wire_ctrl_stage7[102] = counter_w[0]; 
  assign wire_ctrl_stage7[103] = counter_w[0]; 
  assign wire_ctrl_stage7[104] = counter_w[0]; 
  assign wire_ctrl_stage7[105] = counter_w[0]; 
  assign wire_ctrl_stage7[106] = counter_w[0]; 
  assign wire_ctrl_stage7[107] = counter_w[0]; 
  assign wire_ctrl_stage7[108] = counter_w[0]; 
  assign wire_ctrl_stage7[109] = counter_w[0]; 
  assign wire_ctrl_stage7[110] = counter_w[0]; 
  assign wire_ctrl_stage7[111] = counter_w[0]; 
  assign wire_ctrl_stage7[112] = counter_w[0]; 
  assign wire_ctrl_stage7[113] = counter_w[0]; 
  assign wire_ctrl_stage7[114] = counter_w[0]; 
  assign wire_ctrl_stage7[115] = counter_w[0]; 
  assign wire_ctrl_stage7[116] = counter_w[0]; 
  assign wire_ctrl_stage7[117] = counter_w[0]; 
  assign wire_ctrl_stage7[118] = counter_w[0]; 
  assign wire_ctrl_stage7[119] = counter_w[0]; 
  assign wire_ctrl_stage7[120] = counter_w[0]; 
  assign wire_ctrl_stage7[121] = counter_w[0]; 
  assign wire_ctrl_stage7[122] = counter_w[0]; 
  assign wire_ctrl_stage7[123] = counter_w[0]; 
  assign wire_ctrl_stage7[124] = counter_w[0]; 
  assign wire_ctrl_stage7[125] = counter_w[0]; 
  assign wire_ctrl_stage7[126] = counter_w[0]; 
  assign wire_ctrl_stage7[127] = counter_w[0]; 
  
  assign in_start_stage0 = in_start;    
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = out_start_w;    
  
endmodule                        


module switches_stage_st0_0_R(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
ctrl,                            
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;                   
  input [128-1:0] ctrl;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  switch_2_2 switch_inst_0(.inData_0(wireIn[0]), .inData_1(wireIn[1]), .outData_0(wireOut[0]), .outData_1(wireOut[1]), .ctrl(ctrl[0]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_1(.inData_0(wireIn[2]), .inData_1(wireIn[3]), .outData_0(wireOut[2]), .outData_1(wireOut[3]), .ctrl(ctrl[1]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_2(.inData_0(wireIn[4]), .inData_1(wireIn[5]), .outData_0(wireOut[4]), .outData_1(wireOut[5]), .ctrl(ctrl[2]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_3(.inData_0(wireIn[6]), .inData_1(wireIn[7]), .outData_0(wireOut[6]), .outData_1(wireOut[7]), .ctrl(ctrl[3]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_4(.inData_0(wireIn[8]), .inData_1(wireIn[9]), .outData_0(wireOut[8]), .outData_1(wireOut[9]), .ctrl(ctrl[4]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_5(.inData_0(wireIn[10]), .inData_1(wireIn[11]), .outData_0(wireOut[10]), .outData_1(wireOut[11]), .ctrl(ctrl[5]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_6(.inData_0(wireIn[12]), .inData_1(wireIn[13]), .outData_0(wireOut[12]), .outData_1(wireOut[13]), .ctrl(ctrl[6]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_7(.inData_0(wireIn[14]), .inData_1(wireIn[15]), .outData_0(wireOut[14]), .outData_1(wireOut[15]), .ctrl(ctrl[7]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_8(.inData_0(wireIn[16]), .inData_1(wireIn[17]), .outData_0(wireOut[16]), .outData_1(wireOut[17]), .ctrl(ctrl[8]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_9(.inData_0(wireIn[18]), .inData_1(wireIn[19]), .outData_0(wireOut[18]), .outData_1(wireOut[19]), .ctrl(ctrl[9]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_10(.inData_0(wireIn[20]), .inData_1(wireIn[21]), .outData_0(wireOut[20]), .outData_1(wireOut[21]), .ctrl(ctrl[10]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_11(.inData_0(wireIn[22]), .inData_1(wireIn[23]), .outData_0(wireOut[22]), .outData_1(wireOut[23]), .ctrl(ctrl[11]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_12(.inData_0(wireIn[24]), .inData_1(wireIn[25]), .outData_0(wireOut[24]), .outData_1(wireOut[25]), .ctrl(ctrl[12]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_13(.inData_0(wireIn[26]), .inData_1(wireIn[27]), .outData_0(wireOut[26]), .outData_1(wireOut[27]), .ctrl(ctrl[13]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_14(.inData_0(wireIn[28]), .inData_1(wireIn[29]), .outData_0(wireOut[28]), .outData_1(wireOut[29]), .ctrl(ctrl[14]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_15(.inData_0(wireIn[30]), .inData_1(wireIn[31]), .outData_0(wireOut[30]), .outData_1(wireOut[31]), .ctrl(ctrl[15]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_16(.inData_0(wireIn[32]), .inData_1(wireIn[33]), .outData_0(wireOut[32]), .outData_1(wireOut[33]), .ctrl(ctrl[16]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_17(.inData_0(wireIn[34]), .inData_1(wireIn[35]), .outData_0(wireOut[34]), .outData_1(wireOut[35]), .ctrl(ctrl[17]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_18(.inData_0(wireIn[36]), .inData_1(wireIn[37]), .outData_0(wireOut[36]), .outData_1(wireOut[37]), .ctrl(ctrl[18]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_19(.inData_0(wireIn[38]), .inData_1(wireIn[39]), .outData_0(wireOut[38]), .outData_1(wireOut[39]), .ctrl(ctrl[19]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_20(.inData_0(wireIn[40]), .inData_1(wireIn[41]), .outData_0(wireOut[40]), .outData_1(wireOut[41]), .ctrl(ctrl[20]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_21(.inData_0(wireIn[42]), .inData_1(wireIn[43]), .outData_0(wireOut[42]), .outData_1(wireOut[43]), .ctrl(ctrl[21]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_22(.inData_0(wireIn[44]), .inData_1(wireIn[45]), .outData_0(wireOut[44]), .outData_1(wireOut[45]), .ctrl(ctrl[22]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_23(.inData_0(wireIn[46]), .inData_1(wireIn[47]), .outData_0(wireOut[46]), .outData_1(wireOut[47]), .ctrl(ctrl[23]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_24(.inData_0(wireIn[48]), .inData_1(wireIn[49]), .outData_0(wireOut[48]), .outData_1(wireOut[49]), .ctrl(ctrl[24]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_25(.inData_0(wireIn[50]), .inData_1(wireIn[51]), .outData_0(wireOut[50]), .outData_1(wireOut[51]), .ctrl(ctrl[25]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_26(.inData_0(wireIn[52]), .inData_1(wireIn[53]), .outData_0(wireOut[52]), .outData_1(wireOut[53]), .ctrl(ctrl[26]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_27(.inData_0(wireIn[54]), .inData_1(wireIn[55]), .outData_0(wireOut[54]), .outData_1(wireOut[55]), .ctrl(ctrl[27]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_28(.inData_0(wireIn[56]), .inData_1(wireIn[57]), .outData_0(wireOut[56]), .outData_1(wireOut[57]), .ctrl(ctrl[28]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_29(.inData_0(wireIn[58]), .inData_1(wireIn[59]), .outData_0(wireOut[58]), .outData_1(wireOut[59]), .ctrl(ctrl[29]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_30(.inData_0(wireIn[60]), .inData_1(wireIn[61]), .outData_0(wireOut[60]), .outData_1(wireOut[61]), .ctrl(ctrl[30]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_31(.inData_0(wireIn[62]), .inData_1(wireIn[63]), .outData_0(wireOut[62]), .outData_1(wireOut[63]), .ctrl(ctrl[31]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_32(.inData_0(wireIn[64]), .inData_1(wireIn[65]), .outData_0(wireOut[64]), .outData_1(wireOut[65]), .ctrl(ctrl[32]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_33(.inData_0(wireIn[66]), .inData_1(wireIn[67]), .outData_0(wireOut[66]), .outData_1(wireOut[67]), .ctrl(ctrl[33]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_34(.inData_0(wireIn[68]), .inData_1(wireIn[69]), .outData_0(wireOut[68]), .outData_1(wireOut[69]), .ctrl(ctrl[34]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_35(.inData_0(wireIn[70]), .inData_1(wireIn[71]), .outData_0(wireOut[70]), .outData_1(wireOut[71]), .ctrl(ctrl[35]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_36(.inData_0(wireIn[72]), .inData_1(wireIn[73]), .outData_0(wireOut[72]), .outData_1(wireOut[73]), .ctrl(ctrl[36]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_37(.inData_0(wireIn[74]), .inData_1(wireIn[75]), .outData_0(wireOut[74]), .outData_1(wireOut[75]), .ctrl(ctrl[37]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_38(.inData_0(wireIn[76]), .inData_1(wireIn[77]), .outData_0(wireOut[76]), .outData_1(wireOut[77]), .ctrl(ctrl[38]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_39(.inData_0(wireIn[78]), .inData_1(wireIn[79]), .outData_0(wireOut[78]), .outData_1(wireOut[79]), .ctrl(ctrl[39]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_40(.inData_0(wireIn[80]), .inData_1(wireIn[81]), .outData_0(wireOut[80]), .outData_1(wireOut[81]), .ctrl(ctrl[40]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_41(.inData_0(wireIn[82]), .inData_1(wireIn[83]), .outData_0(wireOut[82]), .outData_1(wireOut[83]), .ctrl(ctrl[41]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_42(.inData_0(wireIn[84]), .inData_1(wireIn[85]), .outData_0(wireOut[84]), .outData_1(wireOut[85]), .ctrl(ctrl[42]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_43(.inData_0(wireIn[86]), .inData_1(wireIn[87]), .outData_0(wireOut[86]), .outData_1(wireOut[87]), .ctrl(ctrl[43]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_44(.inData_0(wireIn[88]), .inData_1(wireIn[89]), .outData_0(wireOut[88]), .outData_1(wireOut[89]), .ctrl(ctrl[44]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_45(.inData_0(wireIn[90]), .inData_1(wireIn[91]), .outData_0(wireOut[90]), .outData_1(wireOut[91]), .ctrl(ctrl[45]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_46(.inData_0(wireIn[92]), .inData_1(wireIn[93]), .outData_0(wireOut[92]), .outData_1(wireOut[93]), .ctrl(ctrl[46]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_47(.inData_0(wireIn[94]), .inData_1(wireIn[95]), .outData_0(wireOut[94]), .outData_1(wireOut[95]), .ctrl(ctrl[47]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_48(.inData_0(wireIn[96]), .inData_1(wireIn[97]), .outData_0(wireOut[96]), .outData_1(wireOut[97]), .ctrl(ctrl[48]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_49(.inData_0(wireIn[98]), .inData_1(wireIn[99]), .outData_0(wireOut[98]), .outData_1(wireOut[99]), .ctrl(ctrl[49]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_50(.inData_0(wireIn[100]), .inData_1(wireIn[101]), .outData_0(wireOut[100]), .outData_1(wireOut[101]), .ctrl(ctrl[50]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_51(.inData_0(wireIn[102]), .inData_1(wireIn[103]), .outData_0(wireOut[102]), .outData_1(wireOut[103]), .ctrl(ctrl[51]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_52(.inData_0(wireIn[104]), .inData_1(wireIn[105]), .outData_0(wireOut[104]), .outData_1(wireOut[105]), .ctrl(ctrl[52]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_53(.inData_0(wireIn[106]), .inData_1(wireIn[107]), .outData_0(wireOut[106]), .outData_1(wireOut[107]), .ctrl(ctrl[53]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_54(.inData_0(wireIn[108]), .inData_1(wireIn[109]), .outData_0(wireOut[108]), .outData_1(wireOut[109]), .ctrl(ctrl[54]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_55(.inData_0(wireIn[110]), .inData_1(wireIn[111]), .outData_0(wireOut[110]), .outData_1(wireOut[111]), .ctrl(ctrl[55]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_56(.inData_0(wireIn[112]), .inData_1(wireIn[113]), .outData_0(wireOut[112]), .outData_1(wireOut[113]), .ctrl(ctrl[56]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_57(.inData_0(wireIn[114]), .inData_1(wireIn[115]), .outData_0(wireOut[114]), .outData_1(wireOut[115]), .ctrl(ctrl[57]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_58(.inData_0(wireIn[116]), .inData_1(wireIn[117]), .outData_0(wireOut[116]), .outData_1(wireOut[117]), .ctrl(ctrl[58]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_59(.inData_0(wireIn[118]), .inData_1(wireIn[119]), .outData_0(wireOut[118]), .outData_1(wireOut[119]), .ctrl(ctrl[59]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_60(.inData_0(wireIn[120]), .inData_1(wireIn[121]), .outData_0(wireOut[120]), .outData_1(wireOut[121]), .ctrl(ctrl[60]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_61(.inData_0(wireIn[122]), .inData_1(wireIn[123]), .outData_0(wireOut[122]), .outData_1(wireOut[123]), .ctrl(ctrl[61]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_62(.inData_0(wireIn[124]), .inData_1(wireIn[125]), .outData_0(wireOut[124]), .outData_1(wireOut[125]), .ctrl(ctrl[62]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_63(.inData_0(wireIn[126]), .inData_1(wireIn[127]), .outData_0(wireOut[126]), .outData_1(wireOut[127]), .ctrl(ctrl[63]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_64(.inData_0(wireIn[128]), .inData_1(wireIn[129]), .outData_0(wireOut[128]), .outData_1(wireOut[129]), .ctrl(ctrl[64]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_65(.inData_0(wireIn[130]), .inData_1(wireIn[131]), .outData_0(wireOut[130]), .outData_1(wireOut[131]), .ctrl(ctrl[65]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_66(.inData_0(wireIn[132]), .inData_1(wireIn[133]), .outData_0(wireOut[132]), .outData_1(wireOut[133]), .ctrl(ctrl[66]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_67(.inData_0(wireIn[134]), .inData_1(wireIn[135]), .outData_0(wireOut[134]), .outData_1(wireOut[135]), .ctrl(ctrl[67]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_68(.inData_0(wireIn[136]), .inData_1(wireIn[137]), .outData_0(wireOut[136]), .outData_1(wireOut[137]), .ctrl(ctrl[68]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_69(.inData_0(wireIn[138]), .inData_1(wireIn[139]), .outData_0(wireOut[138]), .outData_1(wireOut[139]), .ctrl(ctrl[69]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_70(.inData_0(wireIn[140]), .inData_1(wireIn[141]), .outData_0(wireOut[140]), .outData_1(wireOut[141]), .ctrl(ctrl[70]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_71(.inData_0(wireIn[142]), .inData_1(wireIn[143]), .outData_0(wireOut[142]), .outData_1(wireOut[143]), .ctrl(ctrl[71]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_72(.inData_0(wireIn[144]), .inData_1(wireIn[145]), .outData_0(wireOut[144]), .outData_1(wireOut[145]), .ctrl(ctrl[72]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_73(.inData_0(wireIn[146]), .inData_1(wireIn[147]), .outData_0(wireOut[146]), .outData_1(wireOut[147]), .ctrl(ctrl[73]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_74(.inData_0(wireIn[148]), .inData_1(wireIn[149]), .outData_0(wireOut[148]), .outData_1(wireOut[149]), .ctrl(ctrl[74]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_75(.inData_0(wireIn[150]), .inData_1(wireIn[151]), .outData_0(wireOut[150]), .outData_1(wireOut[151]), .ctrl(ctrl[75]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_76(.inData_0(wireIn[152]), .inData_1(wireIn[153]), .outData_0(wireOut[152]), .outData_1(wireOut[153]), .ctrl(ctrl[76]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_77(.inData_0(wireIn[154]), .inData_1(wireIn[155]), .outData_0(wireOut[154]), .outData_1(wireOut[155]), .ctrl(ctrl[77]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_78(.inData_0(wireIn[156]), .inData_1(wireIn[157]), .outData_0(wireOut[156]), .outData_1(wireOut[157]), .ctrl(ctrl[78]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_79(.inData_0(wireIn[158]), .inData_1(wireIn[159]), .outData_0(wireOut[158]), .outData_1(wireOut[159]), .ctrl(ctrl[79]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_80(.inData_0(wireIn[160]), .inData_1(wireIn[161]), .outData_0(wireOut[160]), .outData_1(wireOut[161]), .ctrl(ctrl[80]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_81(.inData_0(wireIn[162]), .inData_1(wireIn[163]), .outData_0(wireOut[162]), .outData_1(wireOut[163]), .ctrl(ctrl[81]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_82(.inData_0(wireIn[164]), .inData_1(wireIn[165]), .outData_0(wireOut[164]), .outData_1(wireOut[165]), .ctrl(ctrl[82]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_83(.inData_0(wireIn[166]), .inData_1(wireIn[167]), .outData_0(wireOut[166]), .outData_1(wireOut[167]), .ctrl(ctrl[83]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_84(.inData_0(wireIn[168]), .inData_1(wireIn[169]), .outData_0(wireOut[168]), .outData_1(wireOut[169]), .ctrl(ctrl[84]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_85(.inData_0(wireIn[170]), .inData_1(wireIn[171]), .outData_0(wireOut[170]), .outData_1(wireOut[171]), .ctrl(ctrl[85]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_86(.inData_0(wireIn[172]), .inData_1(wireIn[173]), .outData_0(wireOut[172]), .outData_1(wireOut[173]), .ctrl(ctrl[86]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_87(.inData_0(wireIn[174]), .inData_1(wireIn[175]), .outData_0(wireOut[174]), .outData_1(wireOut[175]), .ctrl(ctrl[87]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_88(.inData_0(wireIn[176]), .inData_1(wireIn[177]), .outData_0(wireOut[176]), .outData_1(wireOut[177]), .ctrl(ctrl[88]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_89(.inData_0(wireIn[178]), .inData_1(wireIn[179]), .outData_0(wireOut[178]), .outData_1(wireOut[179]), .ctrl(ctrl[89]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_90(.inData_0(wireIn[180]), .inData_1(wireIn[181]), .outData_0(wireOut[180]), .outData_1(wireOut[181]), .ctrl(ctrl[90]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_91(.inData_0(wireIn[182]), .inData_1(wireIn[183]), .outData_0(wireOut[182]), .outData_1(wireOut[183]), .ctrl(ctrl[91]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_92(.inData_0(wireIn[184]), .inData_1(wireIn[185]), .outData_0(wireOut[184]), .outData_1(wireOut[185]), .ctrl(ctrl[92]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_93(.inData_0(wireIn[186]), .inData_1(wireIn[187]), .outData_0(wireOut[186]), .outData_1(wireOut[187]), .ctrl(ctrl[93]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_94(.inData_0(wireIn[188]), .inData_1(wireIn[189]), .outData_0(wireOut[188]), .outData_1(wireOut[189]), .ctrl(ctrl[94]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_95(.inData_0(wireIn[190]), .inData_1(wireIn[191]), .outData_0(wireOut[190]), .outData_1(wireOut[191]), .ctrl(ctrl[95]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_96(.inData_0(wireIn[192]), .inData_1(wireIn[193]), .outData_0(wireOut[192]), .outData_1(wireOut[193]), .ctrl(ctrl[96]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_97(.inData_0(wireIn[194]), .inData_1(wireIn[195]), .outData_0(wireOut[194]), .outData_1(wireOut[195]), .ctrl(ctrl[97]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_98(.inData_0(wireIn[196]), .inData_1(wireIn[197]), .outData_0(wireOut[196]), .outData_1(wireOut[197]), .ctrl(ctrl[98]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_99(.inData_0(wireIn[198]), .inData_1(wireIn[199]), .outData_0(wireOut[198]), .outData_1(wireOut[199]), .ctrl(ctrl[99]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_100(.inData_0(wireIn[200]), .inData_1(wireIn[201]), .outData_0(wireOut[200]), .outData_1(wireOut[201]), .ctrl(ctrl[100]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_101(.inData_0(wireIn[202]), .inData_1(wireIn[203]), .outData_0(wireOut[202]), .outData_1(wireOut[203]), .ctrl(ctrl[101]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_102(.inData_0(wireIn[204]), .inData_1(wireIn[205]), .outData_0(wireOut[204]), .outData_1(wireOut[205]), .ctrl(ctrl[102]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_103(.inData_0(wireIn[206]), .inData_1(wireIn[207]), .outData_0(wireOut[206]), .outData_1(wireOut[207]), .ctrl(ctrl[103]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_104(.inData_0(wireIn[208]), .inData_1(wireIn[209]), .outData_0(wireOut[208]), .outData_1(wireOut[209]), .ctrl(ctrl[104]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_105(.inData_0(wireIn[210]), .inData_1(wireIn[211]), .outData_0(wireOut[210]), .outData_1(wireOut[211]), .ctrl(ctrl[105]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_106(.inData_0(wireIn[212]), .inData_1(wireIn[213]), .outData_0(wireOut[212]), .outData_1(wireOut[213]), .ctrl(ctrl[106]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_107(.inData_0(wireIn[214]), .inData_1(wireIn[215]), .outData_0(wireOut[214]), .outData_1(wireOut[215]), .ctrl(ctrl[107]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_108(.inData_0(wireIn[216]), .inData_1(wireIn[217]), .outData_0(wireOut[216]), .outData_1(wireOut[217]), .ctrl(ctrl[108]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_109(.inData_0(wireIn[218]), .inData_1(wireIn[219]), .outData_0(wireOut[218]), .outData_1(wireOut[219]), .ctrl(ctrl[109]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_110(.inData_0(wireIn[220]), .inData_1(wireIn[221]), .outData_0(wireOut[220]), .outData_1(wireOut[221]), .ctrl(ctrl[110]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_111(.inData_0(wireIn[222]), .inData_1(wireIn[223]), .outData_0(wireOut[222]), .outData_1(wireOut[223]), .ctrl(ctrl[111]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_112(.inData_0(wireIn[224]), .inData_1(wireIn[225]), .outData_0(wireOut[224]), .outData_1(wireOut[225]), .ctrl(ctrl[112]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_113(.inData_0(wireIn[226]), .inData_1(wireIn[227]), .outData_0(wireOut[226]), .outData_1(wireOut[227]), .ctrl(ctrl[113]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_114(.inData_0(wireIn[228]), .inData_1(wireIn[229]), .outData_0(wireOut[228]), .outData_1(wireOut[229]), .ctrl(ctrl[114]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_115(.inData_0(wireIn[230]), .inData_1(wireIn[231]), .outData_0(wireOut[230]), .outData_1(wireOut[231]), .ctrl(ctrl[115]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_116(.inData_0(wireIn[232]), .inData_1(wireIn[233]), .outData_0(wireOut[232]), .outData_1(wireOut[233]), .ctrl(ctrl[116]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_117(.inData_0(wireIn[234]), .inData_1(wireIn[235]), .outData_0(wireOut[234]), .outData_1(wireOut[235]), .ctrl(ctrl[117]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_118(.inData_0(wireIn[236]), .inData_1(wireIn[237]), .outData_0(wireOut[236]), .outData_1(wireOut[237]), .ctrl(ctrl[118]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_119(.inData_0(wireIn[238]), .inData_1(wireIn[239]), .outData_0(wireOut[238]), .outData_1(wireOut[239]), .ctrl(ctrl[119]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_120(.inData_0(wireIn[240]), .inData_1(wireIn[241]), .outData_0(wireOut[240]), .outData_1(wireOut[241]), .ctrl(ctrl[120]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_121(.inData_0(wireIn[242]), .inData_1(wireIn[243]), .outData_0(wireOut[242]), .outData_1(wireOut[243]), .ctrl(ctrl[121]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_122(.inData_0(wireIn[244]), .inData_1(wireIn[245]), .outData_0(wireOut[244]), .outData_1(wireOut[245]), .ctrl(ctrl[122]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_123(.inData_0(wireIn[246]), .inData_1(wireIn[247]), .outData_0(wireOut[246]), .outData_1(wireOut[247]), .ctrl(ctrl[123]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_124(.inData_0(wireIn[248]), .inData_1(wireIn[249]), .outData_0(wireOut[248]), .outData_1(wireOut[249]), .ctrl(ctrl[124]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_125(.inData_0(wireIn[250]), .inData_1(wireIn[251]), .outData_0(wireOut[250]), .outData_1(wireOut[251]), .ctrl(ctrl[125]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_126(.inData_0(wireIn[252]), .inData_1(wireIn[253]), .outData_0(wireOut[252]), .outData_1(wireOut[253]), .ctrl(ctrl[126]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_127(.inData_0(wireIn[254]), .inData_1(wireIn[255]), .outData_0(wireOut[254]), .outData_1(wireOut[255]), .ctrl(ctrl[127]), .clk(clk), .rst(rst));
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module wireCon_dp256_st0_R(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  assign wireOut[0] = wireIn[0];    
  assign wireOut[1] = wireIn[128];    
  assign wireOut[2] = wireIn[1];    
  assign wireOut[3] = wireIn[129];    
  assign wireOut[4] = wireIn[2];    
  assign wireOut[5] = wireIn[130];    
  assign wireOut[6] = wireIn[3];    
  assign wireOut[7] = wireIn[131];    
  assign wireOut[8] = wireIn[4];    
  assign wireOut[9] = wireIn[132];    
  assign wireOut[10] = wireIn[5];    
  assign wireOut[11] = wireIn[133];    
  assign wireOut[12] = wireIn[6];    
  assign wireOut[13] = wireIn[134];    
  assign wireOut[14] = wireIn[7];    
  assign wireOut[15] = wireIn[135];    
  assign wireOut[16] = wireIn[8];    
  assign wireOut[17] = wireIn[136];    
  assign wireOut[18] = wireIn[9];    
  assign wireOut[19] = wireIn[137];    
  assign wireOut[20] = wireIn[10];    
  assign wireOut[21] = wireIn[138];    
  assign wireOut[22] = wireIn[11];    
  assign wireOut[23] = wireIn[139];    
  assign wireOut[24] = wireIn[12];    
  assign wireOut[25] = wireIn[140];    
  assign wireOut[26] = wireIn[13];    
  assign wireOut[27] = wireIn[141];    
  assign wireOut[28] = wireIn[14];    
  assign wireOut[29] = wireIn[142];    
  assign wireOut[30] = wireIn[15];    
  assign wireOut[31] = wireIn[143];    
  assign wireOut[32] = wireIn[16];    
  assign wireOut[33] = wireIn[144];    
  assign wireOut[34] = wireIn[17];    
  assign wireOut[35] = wireIn[145];    
  assign wireOut[36] = wireIn[18];    
  assign wireOut[37] = wireIn[146];    
  assign wireOut[38] = wireIn[19];    
  assign wireOut[39] = wireIn[147];    
  assign wireOut[40] = wireIn[20];    
  assign wireOut[41] = wireIn[148];    
  assign wireOut[42] = wireIn[21];    
  assign wireOut[43] = wireIn[149];    
  assign wireOut[44] = wireIn[22];    
  assign wireOut[45] = wireIn[150];    
  assign wireOut[46] = wireIn[23];    
  assign wireOut[47] = wireIn[151];    
  assign wireOut[48] = wireIn[24];    
  assign wireOut[49] = wireIn[152];    
  assign wireOut[50] = wireIn[25];    
  assign wireOut[51] = wireIn[153];    
  assign wireOut[52] = wireIn[26];    
  assign wireOut[53] = wireIn[154];    
  assign wireOut[54] = wireIn[27];    
  assign wireOut[55] = wireIn[155];    
  assign wireOut[56] = wireIn[28];    
  assign wireOut[57] = wireIn[156];    
  assign wireOut[58] = wireIn[29];    
  assign wireOut[59] = wireIn[157];    
  assign wireOut[60] = wireIn[30];    
  assign wireOut[61] = wireIn[158];    
  assign wireOut[62] = wireIn[31];    
  assign wireOut[63] = wireIn[159];    
  assign wireOut[64] = wireIn[32];    
  assign wireOut[65] = wireIn[160];    
  assign wireOut[66] = wireIn[33];    
  assign wireOut[67] = wireIn[161];    
  assign wireOut[68] = wireIn[34];    
  assign wireOut[69] = wireIn[162];    
  assign wireOut[70] = wireIn[35];    
  assign wireOut[71] = wireIn[163];    
  assign wireOut[72] = wireIn[36];    
  assign wireOut[73] = wireIn[164];    
  assign wireOut[74] = wireIn[37];    
  assign wireOut[75] = wireIn[165];    
  assign wireOut[76] = wireIn[38];    
  assign wireOut[77] = wireIn[166];    
  assign wireOut[78] = wireIn[39];    
  assign wireOut[79] = wireIn[167];    
  assign wireOut[80] = wireIn[40];    
  assign wireOut[81] = wireIn[168];    
  assign wireOut[82] = wireIn[41];    
  assign wireOut[83] = wireIn[169];    
  assign wireOut[84] = wireIn[42];    
  assign wireOut[85] = wireIn[170];    
  assign wireOut[86] = wireIn[43];    
  assign wireOut[87] = wireIn[171];    
  assign wireOut[88] = wireIn[44];    
  assign wireOut[89] = wireIn[172];    
  assign wireOut[90] = wireIn[45];    
  assign wireOut[91] = wireIn[173];    
  assign wireOut[92] = wireIn[46];    
  assign wireOut[93] = wireIn[174];    
  assign wireOut[94] = wireIn[47];    
  assign wireOut[95] = wireIn[175];    
  assign wireOut[96] = wireIn[48];    
  assign wireOut[97] = wireIn[176];    
  assign wireOut[98] = wireIn[49];    
  assign wireOut[99] = wireIn[177];    
  assign wireOut[100] = wireIn[50];    
  assign wireOut[101] = wireIn[178];    
  assign wireOut[102] = wireIn[51];    
  assign wireOut[103] = wireIn[179];    
  assign wireOut[104] = wireIn[52];    
  assign wireOut[105] = wireIn[180];    
  assign wireOut[106] = wireIn[53];    
  assign wireOut[107] = wireIn[181];    
  assign wireOut[108] = wireIn[54];    
  assign wireOut[109] = wireIn[182];    
  assign wireOut[110] = wireIn[55];    
  assign wireOut[111] = wireIn[183];    
  assign wireOut[112] = wireIn[56];    
  assign wireOut[113] = wireIn[184];    
  assign wireOut[114] = wireIn[57];    
  assign wireOut[115] = wireIn[185];    
  assign wireOut[116] = wireIn[58];    
  assign wireOut[117] = wireIn[186];    
  assign wireOut[118] = wireIn[59];    
  assign wireOut[119] = wireIn[187];    
  assign wireOut[120] = wireIn[60];    
  assign wireOut[121] = wireIn[188];    
  assign wireOut[122] = wireIn[61];    
  assign wireOut[123] = wireIn[189];    
  assign wireOut[124] = wireIn[62];    
  assign wireOut[125] = wireIn[190];    
  assign wireOut[126] = wireIn[63];    
  assign wireOut[127] = wireIn[191];    
  assign wireOut[128] = wireIn[64];    
  assign wireOut[129] = wireIn[192];    
  assign wireOut[130] = wireIn[65];    
  assign wireOut[131] = wireIn[193];    
  assign wireOut[132] = wireIn[66];    
  assign wireOut[133] = wireIn[194];    
  assign wireOut[134] = wireIn[67];    
  assign wireOut[135] = wireIn[195];    
  assign wireOut[136] = wireIn[68];    
  assign wireOut[137] = wireIn[196];    
  assign wireOut[138] = wireIn[69];    
  assign wireOut[139] = wireIn[197];    
  assign wireOut[140] = wireIn[70];    
  assign wireOut[141] = wireIn[198];    
  assign wireOut[142] = wireIn[71];    
  assign wireOut[143] = wireIn[199];    
  assign wireOut[144] = wireIn[72];    
  assign wireOut[145] = wireIn[200];    
  assign wireOut[146] = wireIn[73];    
  assign wireOut[147] = wireIn[201];    
  assign wireOut[148] = wireIn[74];    
  assign wireOut[149] = wireIn[202];    
  assign wireOut[150] = wireIn[75];    
  assign wireOut[151] = wireIn[203];    
  assign wireOut[152] = wireIn[76];    
  assign wireOut[153] = wireIn[204];    
  assign wireOut[154] = wireIn[77];    
  assign wireOut[155] = wireIn[205];    
  assign wireOut[156] = wireIn[78];    
  assign wireOut[157] = wireIn[206];    
  assign wireOut[158] = wireIn[79];    
  assign wireOut[159] = wireIn[207];    
  assign wireOut[160] = wireIn[80];    
  assign wireOut[161] = wireIn[208];    
  assign wireOut[162] = wireIn[81];    
  assign wireOut[163] = wireIn[209];    
  assign wireOut[164] = wireIn[82];    
  assign wireOut[165] = wireIn[210];    
  assign wireOut[166] = wireIn[83];    
  assign wireOut[167] = wireIn[211];    
  assign wireOut[168] = wireIn[84];    
  assign wireOut[169] = wireIn[212];    
  assign wireOut[170] = wireIn[85];    
  assign wireOut[171] = wireIn[213];    
  assign wireOut[172] = wireIn[86];    
  assign wireOut[173] = wireIn[214];    
  assign wireOut[174] = wireIn[87];    
  assign wireOut[175] = wireIn[215];    
  assign wireOut[176] = wireIn[88];    
  assign wireOut[177] = wireIn[216];    
  assign wireOut[178] = wireIn[89];    
  assign wireOut[179] = wireIn[217];    
  assign wireOut[180] = wireIn[90];    
  assign wireOut[181] = wireIn[218];    
  assign wireOut[182] = wireIn[91];    
  assign wireOut[183] = wireIn[219];    
  assign wireOut[184] = wireIn[92];    
  assign wireOut[185] = wireIn[220];    
  assign wireOut[186] = wireIn[93];    
  assign wireOut[187] = wireIn[221];    
  assign wireOut[188] = wireIn[94];    
  assign wireOut[189] = wireIn[222];    
  assign wireOut[190] = wireIn[95];    
  assign wireOut[191] = wireIn[223];    
  assign wireOut[192] = wireIn[96];    
  assign wireOut[193] = wireIn[224];    
  assign wireOut[194] = wireIn[97];    
  assign wireOut[195] = wireIn[225];    
  assign wireOut[196] = wireIn[98];    
  assign wireOut[197] = wireIn[226];    
  assign wireOut[198] = wireIn[99];    
  assign wireOut[199] = wireIn[227];    
  assign wireOut[200] = wireIn[100];    
  assign wireOut[201] = wireIn[228];    
  assign wireOut[202] = wireIn[101];    
  assign wireOut[203] = wireIn[229];    
  assign wireOut[204] = wireIn[102];    
  assign wireOut[205] = wireIn[230];    
  assign wireOut[206] = wireIn[103];    
  assign wireOut[207] = wireIn[231];    
  assign wireOut[208] = wireIn[104];    
  assign wireOut[209] = wireIn[232];    
  assign wireOut[210] = wireIn[105];    
  assign wireOut[211] = wireIn[233];    
  assign wireOut[212] = wireIn[106];    
  assign wireOut[213] = wireIn[234];    
  assign wireOut[214] = wireIn[107];    
  assign wireOut[215] = wireIn[235];    
  assign wireOut[216] = wireIn[108];    
  assign wireOut[217] = wireIn[236];    
  assign wireOut[218] = wireIn[109];    
  assign wireOut[219] = wireIn[237];    
  assign wireOut[220] = wireIn[110];    
  assign wireOut[221] = wireIn[238];    
  assign wireOut[222] = wireIn[111];    
  assign wireOut[223] = wireIn[239];    
  assign wireOut[224] = wireIn[112];    
  assign wireOut[225] = wireIn[240];    
  assign wireOut[226] = wireIn[113];    
  assign wireOut[227] = wireIn[241];    
  assign wireOut[228] = wireIn[114];    
  assign wireOut[229] = wireIn[242];    
  assign wireOut[230] = wireIn[115];    
  assign wireOut[231] = wireIn[243];    
  assign wireOut[232] = wireIn[116];    
  assign wireOut[233] = wireIn[244];    
  assign wireOut[234] = wireIn[117];    
  assign wireOut[235] = wireIn[245];    
  assign wireOut[236] = wireIn[118];    
  assign wireOut[237] = wireIn[246];    
  assign wireOut[238] = wireIn[119];    
  assign wireOut[239] = wireIn[247];    
  assign wireOut[240] = wireIn[120];    
  assign wireOut[241] = wireIn[248];    
  assign wireOut[242] = wireIn[121];    
  assign wireOut[243] = wireIn[249];    
  assign wireOut[244] = wireIn[122];    
  assign wireOut[245] = wireIn[250];    
  assign wireOut[246] = wireIn[123];    
  assign wireOut[247] = wireIn[251];    
  assign wireOut[248] = wireIn[124];    
  assign wireOut[249] = wireIn[252];    
  assign wireOut[250] = wireIn[125];    
  assign wireOut[251] = wireIn[253];    
  assign wireOut[252] = wireIn[126];    
  assign wireOut[253] = wireIn[254];    
  assign wireOut[254] = wireIn[127];    
  assign wireOut[255] = wireIn[255];    
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module switches_stage_st1_0_R(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
ctrl,                            
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;                   
  input [128-1:0] ctrl;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  switch_2_2 switch_inst_0(.inData_0(wireIn[0]), .inData_1(wireIn[1]), .outData_0(wireOut[0]), .outData_1(wireOut[1]), .ctrl(ctrl[0]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_1(.inData_0(wireIn[2]), .inData_1(wireIn[3]), .outData_0(wireOut[2]), .outData_1(wireOut[3]), .ctrl(ctrl[1]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_2(.inData_0(wireIn[4]), .inData_1(wireIn[5]), .outData_0(wireOut[4]), .outData_1(wireOut[5]), .ctrl(ctrl[2]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_3(.inData_0(wireIn[6]), .inData_1(wireIn[7]), .outData_0(wireOut[6]), .outData_1(wireOut[7]), .ctrl(ctrl[3]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_4(.inData_0(wireIn[8]), .inData_1(wireIn[9]), .outData_0(wireOut[8]), .outData_1(wireOut[9]), .ctrl(ctrl[4]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_5(.inData_0(wireIn[10]), .inData_1(wireIn[11]), .outData_0(wireOut[10]), .outData_1(wireOut[11]), .ctrl(ctrl[5]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_6(.inData_0(wireIn[12]), .inData_1(wireIn[13]), .outData_0(wireOut[12]), .outData_1(wireOut[13]), .ctrl(ctrl[6]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_7(.inData_0(wireIn[14]), .inData_1(wireIn[15]), .outData_0(wireOut[14]), .outData_1(wireOut[15]), .ctrl(ctrl[7]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_8(.inData_0(wireIn[16]), .inData_1(wireIn[17]), .outData_0(wireOut[16]), .outData_1(wireOut[17]), .ctrl(ctrl[8]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_9(.inData_0(wireIn[18]), .inData_1(wireIn[19]), .outData_0(wireOut[18]), .outData_1(wireOut[19]), .ctrl(ctrl[9]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_10(.inData_0(wireIn[20]), .inData_1(wireIn[21]), .outData_0(wireOut[20]), .outData_1(wireOut[21]), .ctrl(ctrl[10]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_11(.inData_0(wireIn[22]), .inData_1(wireIn[23]), .outData_0(wireOut[22]), .outData_1(wireOut[23]), .ctrl(ctrl[11]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_12(.inData_0(wireIn[24]), .inData_1(wireIn[25]), .outData_0(wireOut[24]), .outData_1(wireOut[25]), .ctrl(ctrl[12]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_13(.inData_0(wireIn[26]), .inData_1(wireIn[27]), .outData_0(wireOut[26]), .outData_1(wireOut[27]), .ctrl(ctrl[13]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_14(.inData_0(wireIn[28]), .inData_1(wireIn[29]), .outData_0(wireOut[28]), .outData_1(wireOut[29]), .ctrl(ctrl[14]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_15(.inData_0(wireIn[30]), .inData_1(wireIn[31]), .outData_0(wireOut[30]), .outData_1(wireOut[31]), .ctrl(ctrl[15]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_16(.inData_0(wireIn[32]), .inData_1(wireIn[33]), .outData_0(wireOut[32]), .outData_1(wireOut[33]), .ctrl(ctrl[16]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_17(.inData_0(wireIn[34]), .inData_1(wireIn[35]), .outData_0(wireOut[34]), .outData_1(wireOut[35]), .ctrl(ctrl[17]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_18(.inData_0(wireIn[36]), .inData_1(wireIn[37]), .outData_0(wireOut[36]), .outData_1(wireOut[37]), .ctrl(ctrl[18]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_19(.inData_0(wireIn[38]), .inData_1(wireIn[39]), .outData_0(wireOut[38]), .outData_1(wireOut[39]), .ctrl(ctrl[19]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_20(.inData_0(wireIn[40]), .inData_1(wireIn[41]), .outData_0(wireOut[40]), .outData_1(wireOut[41]), .ctrl(ctrl[20]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_21(.inData_0(wireIn[42]), .inData_1(wireIn[43]), .outData_0(wireOut[42]), .outData_1(wireOut[43]), .ctrl(ctrl[21]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_22(.inData_0(wireIn[44]), .inData_1(wireIn[45]), .outData_0(wireOut[44]), .outData_1(wireOut[45]), .ctrl(ctrl[22]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_23(.inData_0(wireIn[46]), .inData_1(wireIn[47]), .outData_0(wireOut[46]), .outData_1(wireOut[47]), .ctrl(ctrl[23]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_24(.inData_0(wireIn[48]), .inData_1(wireIn[49]), .outData_0(wireOut[48]), .outData_1(wireOut[49]), .ctrl(ctrl[24]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_25(.inData_0(wireIn[50]), .inData_1(wireIn[51]), .outData_0(wireOut[50]), .outData_1(wireOut[51]), .ctrl(ctrl[25]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_26(.inData_0(wireIn[52]), .inData_1(wireIn[53]), .outData_0(wireOut[52]), .outData_1(wireOut[53]), .ctrl(ctrl[26]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_27(.inData_0(wireIn[54]), .inData_1(wireIn[55]), .outData_0(wireOut[54]), .outData_1(wireOut[55]), .ctrl(ctrl[27]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_28(.inData_0(wireIn[56]), .inData_1(wireIn[57]), .outData_0(wireOut[56]), .outData_1(wireOut[57]), .ctrl(ctrl[28]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_29(.inData_0(wireIn[58]), .inData_1(wireIn[59]), .outData_0(wireOut[58]), .outData_1(wireOut[59]), .ctrl(ctrl[29]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_30(.inData_0(wireIn[60]), .inData_1(wireIn[61]), .outData_0(wireOut[60]), .outData_1(wireOut[61]), .ctrl(ctrl[30]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_31(.inData_0(wireIn[62]), .inData_1(wireIn[63]), .outData_0(wireOut[62]), .outData_1(wireOut[63]), .ctrl(ctrl[31]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_32(.inData_0(wireIn[64]), .inData_1(wireIn[65]), .outData_0(wireOut[64]), .outData_1(wireOut[65]), .ctrl(ctrl[32]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_33(.inData_0(wireIn[66]), .inData_1(wireIn[67]), .outData_0(wireOut[66]), .outData_1(wireOut[67]), .ctrl(ctrl[33]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_34(.inData_0(wireIn[68]), .inData_1(wireIn[69]), .outData_0(wireOut[68]), .outData_1(wireOut[69]), .ctrl(ctrl[34]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_35(.inData_0(wireIn[70]), .inData_1(wireIn[71]), .outData_0(wireOut[70]), .outData_1(wireOut[71]), .ctrl(ctrl[35]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_36(.inData_0(wireIn[72]), .inData_1(wireIn[73]), .outData_0(wireOut[72]), .outData_1(wireOut[73]), .ctrl(ctrl[36]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_37(.inData_0(wireIn[74]), .inData_1(wireIn[75]), .outData_0(wireOut[74]), .outData_1(wireOut[75]), .ctrl(ctrl[37]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_38(.inData_0(wireIn[76]), .inData_1(wireIn[77]), .outData_0(wireOut[76]), .outData_1(wireOut[77]), .ctrl(ctrl[38]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_39(.inData_0(wireIn[78]), .inData_1(wireIn[79]), .outData_0(wireOut[78]), .outData_1(wireOut[79]), .ctrl(ctrl[39]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_40(.inData_0(wireIn[80]), .inData_1(wireIn[81]), .outData_0(wireOut[80]), .outData_1(wireOut[81]), .ctrl(ctrl[40]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_41(.inData_0(wireIn[82]), .inData_1(wireIn[83]), .outData_0(wireOut[82]), .outData_1(wireOut[83]), .ctrl(ctrl[41]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_42(.inData_0(wireIn[84]), .inData_1(wireIn[85]), .outData_0(wireOut[84]), .outData_1(wireOut[85]), .ctrl(ctrl[42]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_43(.inData_0(wireIn[86]), .inData_1(wireIn[87]), .outData_0(wireOut[86]), .outData_1(wireOut[87]), .ctrl(ctrl[43]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_44(.inData_0(wireIn[88]), .inData_1(wireIn[89]), .outData_0(wireOut[88]), .outData_1(wireOut[89]), .ctrl(ctrl[44]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_45(.inData_0(wireIn[90]), .inData_1(wireIn[91]), .outData_0(wireOut[90]), .outData_1(wireOut[91]), .ctrl(ctrl[45]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_46(.inData_0(wireIn[92]), .inData_1(wireIn[93]), .outData_0(wireOut[92]), .outData_1(wireOut[93]), .ctrl(ctrl[46]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_47(.inData_0(wireIn[94]), .inData_1(wireIn[95]), .outData_0(wireOut[94]), .outData_1(wireOut[95]), .ctrl(ctrl[47]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_48(.inData_0(wireIn[96]), .inData_1(wireIn[97]), .outData_0(wireOut[96]), .outData_1(wireOut[97]), .ctrl(ctrl[48]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_49(.inData_0(wireIn[98]), .inData_1(wireIn[99]), .outData_0(wireOut[98]), .outData_1(wireOut[99]), .ctrl(ctrl[49]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_50(.inData_0(wireIn[100]), .inData_1(wireIn[101]), .outData_0(wireOut[100]), .outData_1(wireOut[101]), .ctrl(ctrl[50]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_51(.inData_0(wireIn[102]), .inData_1(wireIn[103]), .outData_0(wireOut[102]), .outData_1(wireOut[103]), .ctrl(ctrl[51]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_52(.inData_0(wireIn[104]), .inData_1(wireIn[105]), .outData_0(wireOut[104]), .outData_1(wireOut[105]), .ctrl(ctrl[52]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_53(.inData_0(wireIn[106]), .inData_1(wireIn[107]), .outData_0(wireOut[106]), .outData_1(wireOut[107]), .ctrl(ctrl[53]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_54(.inData_0(wireIn[108]), .inData_1(wireIn[109]), .outData_0(wireOut[108]), .outData_1(wireOut[109]), .ctrl(ctrl[54]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_55(.inData_0(wireIn[110]), .inData_1(wireIn[111]), .outData_0(wireOut[110]), .outData_1(wireOut[111]), .ctrl(ctrl[55]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_56(.inData_0(wireIn[112]), .inData_1(wireIn[113]), .outData_0(wireOut[112]), .outData_1(wireOut[113]), .ctrl(ctrl[56]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_57(.inData_0(wireIn[114]), .inData_1(wireIn[115]), .outData_0(wireOut[114]), .outData_1(wireOut[115]), .ctrl(ctrl[57]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_58(.inData_0(wireIn[116]), .inData_1(wireIn[117]), .outData_0(wireOut[116]), .outData_1(wireOut[117]), .ctrl(ctrl[58]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_59(.inData_0(wireIn[118]), .inData_1(wireIn[119]), .outData_0(wireOut[118]), .outData_1(wireOut[119]), .ctrl(ctrl[59]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_60(.inData_0(wireIn[120]), .inData_1(wireIn[121]), .outData_0(wireOut[120]), .outData_1(wireOut[121]), .ctrl(ctrl[60]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_61(.inData_0(wireIn[122]), .inData_1(wireIn[123]), .outData_0(wireOut[122]), .outData_1(wireOut[123]), .ctrl(ctrl[61]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_62(.inData_0(wireIn[124]), .inData_1(wireIn[125]), .outData_0(wireOut[124]), .outData_1(wireOut[125]), .ctrl(ctrl[62]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_63(.inData_0(wireIn[126]), .inData_1(wireIn[127]), .outData_0(wireOut[126]), .outData_1(wireOut[127]), .ctrl(ctrl[63]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_64(.inData_0(wireIn[128]), .inData_1(wireIn[129]), .outData_0(wireOut[128]), .outData_1(wireOut[129]), .ctrl(ctrl[64]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_65(.inData_0(wireIn[130]), .inData_1(wireIn[131]), .outData_0(wireOut[130]), .outData_1(wireOut[131]), .ctrl(ctrl[65]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_66(.inData_0(wireIn[132]), .inData_1(wireIn[133]), .outData_0(wireOut[132]), .outData_1(wireOut[133]), .ctrl(ctrl[66]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_67(.inData_0(wireIn[134]), .inData_1(wireIn[135]), .outData_0(wireOut[134]), .outData_1(wireOut[135]), .ctrl(ctrl[67]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_68(.inData_0(wireIn[136]), .inData_1(wireIn[137]), .outData_0(wireOut[136]), .outData_1(wireOut[137]), .ctrl(ctrl[68]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_69(.inData_0(wireIn[138]), .inData_1(wireIn[139]), .outData_0(wireOut[138]), .outData_1(wireOut[139]), .ctrl(ctrl[69]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_70(.inData_0(wireIn[140]), .inData_1(wireIn[141]), .outData_0(wireOut[140]), .outData_1(wireOut[141]), .ctrl(ctrl[70]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_71(.inData_0(wireIn[142]), .inData_1(wireIn[143]), .outData_0(wireOut[142]), .outData_1(wireOut[143]), .ctrl(ctrl[71]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_72(.inData_0(wireIn[144]), .inData_1(wireIn[145]), .outData_0(wireOut[144]), .outData_1(wireOut[145]), .ctrl(ctrl[72]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_73(.inData_0(wireIn[146]), .inData_1(wireIn[147]), .outData_0(wireOut[146]), .outData_1(wireOut[147]), .ctrl(ctrl[73]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_74(.inData_0(wireIn[148]), .inData_1(wireIn[149]), .outData_0(wireOut[148]), .outData_1(wireOut[149]), .ctrl(ctrl[74]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_75(.inData_0(wireIn[150]), .inData_1(wireIn[151]), .outData_0(wireOut[150]), .outData_1(wireOut[151]), .ctrl(ctrl[75]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_76(.inData_0(wireIn[152]), .inData_1(wireIn[153]), .outData_0(wireOut[152]), .outData_1(wireOut[153]), .ctrl(ctrl[76]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_77(.inData_0(wireIn[154]), .inData_1(wireIn[155]), .outData_0(wireOut[154]), .outData_1(wireOut[155]), .ctrl(ctrl[77]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_78(.inData_0(wireIn[156]), .inData_1(wireIn[157]), .outData_0(wireOut[156]), .outData_1(wireOut[157]), .ctrl(ctrl[78]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_79(.inData_0(wireIn[158]), .inData_1(wireIn[159]), .outData_0(wireOut[158]), .outData_1(wireOut[159]), .ctrl(ctrl[79]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_80(.inData_0(wireIn[160]), .inData_1(wireIn[161]), .outData_0(wireOut[160]), .outData_1(wireOut[161]), .ctrl(ctrl[80]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_81(.inData_0(wireIn[162]), .inData_1(wireIn[163]), .outData_0(wireOut[162]), .outData_1(wireOut[163]), .ctrl(ctrl[81]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_82(.inData_0(wireIn[164]), .inData_1(wireIn[165]), .outData_0(wireOut[164]), .outData_1(wireOut[165]), .ctrl(ctrl[82]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_83(.inData_0(wireIn[166]), .inData_1(wireIn[167]), .outData_0(wireOut[166]), .outData_1(wireOut[167]), .ctrl(ctrl[83]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_84(.inData_0(wireIn[168]), .inData_1(wireIn[169]), .outData_0(wireOut[168]), .outData_1(wireOut[169]), .ctrl(ctrl[84]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_85(.inData_0(wireIn[170]), .inData_1(wireIn[171]), .outData_0(wireOut[170]), .outData_1(wireOut[171]), .ctrl(ctrl[85]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_86(.inData_0(wireIn[172]), .inData_1(wireIn[173]), .outData_0(wireOut[172]), .outData_1(wireOut[173]), .ctrl(ctrl[86]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_87(.inData_0(wireIn[174]), .inData_1(wireIn[175]), .outData_0(wireOut[174]), .outData_1(wireOut[175]), .ctrl(ctrl[87]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_88(.inData_0(wireIn[176]), .inData_1(wireIn[177]), .outData_0(wireOut[176]), .outData_1(wireOut[177]), .ctrl(ctrl[88]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_89(.inData_0(wireIn[178]), .inData_1(wireIn[179]), .outData_0(wireOut[178]), .outData_1(wireOut[179]), .ctrl(ctrl[89]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_90(.inData_0(wireIn[180]), .inData_1(wireIn[181]), .outData_0(wireOut[180]), .outData_1(wireOut[181]), .ctrl(ctrl[90]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_91(.inData_0(wireIn[182]), .inData_1(wireIn[183]), .outData_0(wireOut[182]), .outData_1(wireOut[183]), .ctrl(ctrl[91]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_92(.inData_0(wireIn[184]), .inData_1(wireIn[185]), .outData_0(wireOut[184]), .outData_1(wireOut[185]), .ctrl(ctrl[92]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_93(.inData_0(wireIn[186]), .inData_1(wireIn[187]), .outData_0(wireOut[186]), .outData_1(wireOut[187]), .ctrl(ctrl[93]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_94(.inData_0(wireIn[188]), .inData_1(wireIn[189]), .outData_0(wireOut[188]), .outData_1(wireOut[189]), .ctrl(ctrl[94]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_95(.inData_0(wireIn[190]), .inData_1(wireIn[191]), .outData_0(wireOut[190]), .outData_1(wireOut[191]), .ctrl(ctrl[95]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_96(.inData_0(wireIn[192]), .inData_1(wireIn[193]), .outData_0(wireOut[192]), .outData_1(wireOut[193]), .ctrl(ctrl[96]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_97(.inData_0(wireIn[194]), .inData_1(wireIn[195]), .outData_0(wireOut[194]), .outData_1(wireOut[195]), .ctrl(ctrl[97]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_98(.inData_0(wireIn[196]), .inData_1(wireIn[197]), .outData_0(wireOut[196]), .outData_1(wireOut[197]), .ctrl(ctrl[98]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_99(.inData_0(wireIn[198]), .inData_1(wireIn[199]), .outData_0(wireOut[198]), .outData_1(wireOut[199]), .ctrl(ctrl[99]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_100(.inData_0(wireIn[200]), .inData_1(wireIn[201]), .outData_0(wireOut[200]), .outData_1(wireOut[201]), .ctrl(ctrl[100]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_101(.inData_0(wireIn[202]), .inData_1(wireIn[203]), .outData_0(wireOut[202]), .outData_1(wireOut[203]), .ctrl(ctrl[101]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_102(.inData_0(wireIn[204]), .inData_1(wireIn[205]), .outData_0(wireOut[204]), .outData_1(wireOut[205]), .ctrl(ctrl[102]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_103(.inData_0(wireIn[206]), .inData_1(wireIn[207]), .outData_0(wireOut[206]), .outData_1(wireOut[207]), .ctrl(ctrl[103]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_104(.inData_0(wireIn[208]), .inData_1(wireIn[209]), .outData_0(wireOut[208]), .outData_1(wireOut[209]), .ctrl(ctrl[104]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_105(.inData_0(wireIn[210]), .inData_1(wireIn[211]), .outData_0(wireOut[210]), .outData_1(wireOut[211]), .ctrl(ctrl[105]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_106(.inData_0(wireIn[212]), .inData_1(wireIn[213]), .outData_0(wireOut[212]), .outData_1(wireOut[213]), .ctrl(ctrl[106]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_107(.inData_0(wireIn[214]), .inData_1(wireIn[215]), .outData_0(wireOut[214]), .outData_1(wireOut[215]), .ctrl(ctrl[107]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_108(.inData_0(wireIn[216]), .inData_1(wireIn[217]), .outData_0(wireOut[216]), .outData_1(wireOut[217]), .ctrl(ctrl[108]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_109(.inData_0(wireIn[218]), .inData_1(wireIn[219]), .outData_0(wireOut[218]), .outData_1(wireOut[219]), .ctrl(ctrl[109]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_110(.inData_0(wireIn[220]), .inData_1(wireIn[221]), .outData_0(wireOut[220]), .outData_1(wireOut[221]), .ctrl(ctrl[110]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_111(.inData_0(wireIn[222]), .inData_1(wireIn[223]), .outData_0(wireOut[222]), .outData_1(wireOut[223]), .ctrl(ctrl[111]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_112(.inData_0(wireIn[224]), .inData_1(wireIn[225]), .outData_0(wireOut[224]), .outData_1(wireOut[225]), .ctrl(ctrl[112]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_113(.inData_0(wireIn[226]), .inData_1(wireIn[227]), .outData_0(wireOut[226]), .outData_1(wireOut[227]), .ctrl(ctrl[113]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_114(.inData_0(wireIn[228]), .inData_1(wireIn[229]), .outData_0(wireOut[228]), .outData_1(wireOut[229]), .ctrl(ctrl[114]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_115(.inData_0(wireIn[230]), .inData_1(wireIn[231]), .outData_0(wireOut[230]), .outData_1(wireOut[231]), .ctrl(ctrl[115]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_116(.inData_0(wireIn[232]), .inData_1(wireIn[233]), .outData_0(wireOut[232]), .outData_1(wireOut[233]), .ctrl(ctrl[116]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_117(.inData_0(wireIn[234]), .inData_1(wireIn[235]), .outData_0(wireOut[234]), .outData_1(wireOut[235]), .ctrl(ctrl[117]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_118(.inData_0(wireIn[236]), .inData_1(wireIn[237]), .outData_0(wireOut[236]), .outData_1(wireOut[237]), .ctrl(ctrl[118]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_119(.inData_0(wireIn[238]), .inData_1(wireIn[239]), .outData_0(wireOut[238]), .outData_1(wireOut[239]), .ctrl(ctrl[119]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_120(.inData_0(wireIn[240]), .inData_1(wireIn[241]), .outData_0(wireOut[240]), .outData_1(wireOut[241]), .ctrl(ctrl[120]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_121(.inData_0(wireIn[242]), .inData_1(wireIn[243]), .outData_0(wireOut[242]), .outData_1(wireOut[243]), .ctrl(ctrl[121]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_122(.inData_0(wireIn[244]), .inData_1(wireIn[245]), .outData_0(wireOut[244]), .outData_1(wireOut[245]), .ctrl(ctrl[122]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_123(.inData_0(wireIn[246]), .inData_1(wireIn[247]), .outData_0(wireOut[246]), .outData_1(wireOut[247]), .ctrl(ctrl[123]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_124(.inData_0(wireIn[248]), .inData_1(wireIn[249]), .outData_0(wireOut[248]), .outData_1(wireOut[249]), .ctrl(ctrl[124]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_125(.inData_0(wireIn[250]), .inData_1(wireIn[251]), .outData_0(wireOut[250]), .outData_1(wireOut[251]), .ctrl(ctrl[125]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_126(.inData_0(wireIn[252]), .inData_1(wireIn[253]), .outData_0(wireOut[252]), .outData_1(wireOut[253]), .ctrl(ctrl[126]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_127(.inData_0(wireIn[254]), .inData_1(wireIn[255]), .outData_0(wireOut[254]), .outData_1(wireOut[255]), .ctrl(ctrl[127]), .clk(clk), .rst(rst));
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module wireCon_dp256_st1_R(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  assign wireOut[0] = wireIn[0];    
  assign wireOut[1] = wireIn[64];    
  assign wireOut[2] = wireIn[1];    
  assign wireOut[3] = wireIn[65];    
  assign wireOut[4] = wireIn[2];    
  assign wireOut[5] = wireIn[66];    
  assign wireOut[6] = wireIn[3];    
  assign wireOut[7] = wireIn[67];    
  assign wireOut[8] = wireIn[4];    
  assign wireOut[9] = wireIn[68];    
  assign wireOut[10] = wireIn[5];    
  assign wireOut[11] = wireIn[69];    
  assign wireOut[12] = wireIn[6];    
  assign wireOut[13] = wireIn[70];    
  assign wireOut[14] = wireIn[7];    
  assign wireOut[15] = wireIn[71];    
  assign wireOut[16] = wireIn[8];    
  assign wireOut[17] = wireIn[72];    
  assign wireOut[18] = wireIn[9];    
  assign wireOut[19] = wireIn[73];    
  assign wireOut[20] = wireIn[10];    
  assign wireOut[21] = wireIn[74];    
  assign wireOut[22] = wireIn[11];    
  assign wireOut[23] = wireIn[75];    
  assign wireOut[24] = wireIn[12];    
  assign wireOut[25] = wireIn[76];    
  assign wireOut[26] = wireIn[13];    
  assign wireOut[27] = wireIn[77];    
  assign wireOut[28] = wireIn[14];    
  assign wireOut[29] = wireIn[78];    
  assign wireOut[30] = wireIn[15];    
  assign wireOut[31] = wireIn[79];    
  assign wireOut[32] = wireIn[16];    
  assign wireOut[33] = wireIn[80];    
  assign wireOut[34] = wireIn[17];    
  assign wireOut[35] = wireIn[81];    
  assign wireOut[36] = wireIn[18];    
  assign wireOut[37] = wireIn[82];    
  assign wireOut[38] = wireIn[19];    
  assign wireOut[39] = wireIn[83];    
  assign wireOut[40] = wireIn[20];    
  assign wireOut[41] = wireIn[84];    
  assign wireOut[42] = wireIn[21];    
  assign wireOut[43] = wireIn[85];    
  assign wireOut[44] = wireIn[22];    
  assign wireOut[45] = wireIn[86];    
  assign wireOut[46] = wireIn[23];    
  assign wireOut[47] = wireIn[87];    
  assign wireOut[48] = wireIn[24];    
  assign wireOut[49] = wireIn[88];    
  assign wireOut[50] = wireIn[25];    
  assign wireOut[51] = wireIn[89];    
  assign wireOut[52] = wireIn[26];    
  assign wireOut[53] = wireIn[90];    
  assign wireOut[54] = wireIn[27];    
  assign wireOut[55] = wireIn[91];    
  assign wireOut[56] = wireIn[28];    
  assign wireOut[57] = wireIn[92];    
  assign wireOut[58] = wireIn[29];    
  assign wireOut[59] = wireIn[93];    
  assign wireOut[60] = wireIn[30];    
  assign wireOut[61] = wireIn[94];    
  assign wireOut[62] = wireIn[31];    
  assign wireOut[63] = wireIn[95];    
  assign wireOut[64] = wireIn[32];    
  assign wireOut[65] = wireIn[96];    
  assign wireOut[66] = wireIn[33];    
  assign wireOut[67] = wireIn[97];    
  assign wireOut[68] = wireIn[34];    
  assign wireOut[69] = wireIn[98];    
  assign wireOut[70] = wireIn[35];    
  assign wireOut[71] = wireIn[99];    
  assign wireOut[72] = wireIn[36];    
  assign wireOut[73] = wireIn[100];    
  assign wireOut[74] = wireIn[37];    
  assign wireOut[75] = wireIn[101];    
  assign wireOut[76] = wireIn[38];    
  assign wireOut[77] = wireIn[102];    
  assign wireOut[78] = wireIn[39];    
  assign wireOut[79] = wireIn[103];    
  assign wireOut[80] = wireIn[40];    
  assign wireOut[81] = wireIn[104];    
  assign wireOut[82] = wireIn[41];    
  assign wireOut[83] = wireIn[105];    
  assign wireOut[84] = wireIn[42];    
  assign wireOut[85] = wireIn[106];    
  assign wireOut[86] = wireIn[43];    
  assign wireOut[87] = wireIn[107];    
  assign wireOut[88] = wireIn[44];    
  assign wireOut[89] = wireIn[108];    
  assign wireOut[90] = wireIn[45];    
  assign wireOut[91] = wireIn[109];    
  assign wireOut[92] = wireIn[46];    
  assign wireOut[93] = wireIn[110];    
  assign wireOut[94] = wireIn[47];    
  assign wireOut[95] = wireIn[111];    
  assign wireOut[96] = wireIn[48];    
  assign wireOut[97] = wireIn[112];    
  assign wireOut[98] = wireIn[49];    
  assign wireOut[99] = wireIn[113];    
  assign wireOut[100] = wireIn[50];    
  assign wireOut[101] = wireIn[114];    
  assign wireOut[102] = wireIn[51];    
  assign wireOut[103] = wireIn[115];    
  assign wireOut[104] = wireIn[52];    
  assign wireOut[105] = wireIn[116];    
  assign wireOut[106] = wireIn[53];    
  assign wireOut[107] = wireIn[117];    
  assign wireOut[108] = wireIn[54];    
  assign wireOut[109] = wireIn[118];    
  assign wireOut[110] = wireIn[55];    
  assign wireOut[111] = wireIn[119];    
  assign wireOut[112] = wireIn[56];    
  assign wireOut[113] = wireIn[120];    
  assign wireOut[114] = wireIn[57];    
  assign wireOut[115] = wireIn[121];    
  assign wireOut[116] = wireIn[58];    
  assign wireOut[117] = wireIn[122];    
  assign wireOut[118] = wireIn[59];    
  assign wireOut[119] = wireIn[123];    
  assign wireOut[120] = wireIn[60];    
  assign wireOut[121] = wireIn[124];    
  assign wireOut[122] = wireIn[61];    
  assign wireOut[123] = wireIn[125];    
  assign wireOut[124] = wireIn[62];    
  assign wireOut[125] = wireIn[126];    
  assign wireOut[126] = wireIn[63];    
  assign wireOut[127] = wireIn[127];    
  assign wireOut[128] = wireIn[128];    
  assign wireOut[129] = wireIn[192];    
  assign wireOut[130] = wireIn[129];    
  assign wireOut[131] = wireIn[193];    
  assign wireOut[132] = wireIn[130];    
  assign wireOut[133] = wireIn[194];    
  assign wireOut[134] = wireIn[131];    
  assign wireOut[135] = wireIn[195];    
  assign wireOut[136] = wireIn[132];    
  assign wireOut[137] = wireIn[196];    
  assign wireOut[138] = wireIn[133];    
  assign wireOut[139] = wireIn[197];    
  assign wireOut[140] = wireIn[134];    
  assign wireOut[141] = wireIn[198];    
  assign wireOut[142] = wireIn[135];    
  assign wireOut[143] = wireIn[199];    
  assign wireOut[144] = wireIn[136];    
  assign wireOut[145] = wireIn[200];    
  assign wireOut[146] = wireIn[137];    
  assign wireOut[147] = wireIn[201];    
  assign wireOut[148] = wireIn[138];    
  assign wireOut[149] = wireIn[202];    
  assign wireOut[150] = wireIn[139];    
  assign wireOut[151] = wireIn[203];    
  assign wireOut[152] = wireIn[140];    
  assign wireOut[153] = wireIn[204];    
  assign wireOut[154] = wireIn[141];    
  assign wireOut[155] = wireIn[205];    
  assign wireOut[156] = wireIn[142];    
  assign wireOut[157] = wireIn[206];    
  assign wireOut[158] = wireIn[143];    
  assign wireOut[159] = wireIn[207];    
  assign wireOut[160] = wireIn[144];    
  assign wireOut[161] = wireIn[208];    
  assign wireOut[162] = wireIn[145];    
  assign wireOut[163] = wireIn[209];    
  assign wireOut[164] = wireIn[146];    
  assign wireOut[165] = wireIn[210];    
  assign wireOut[166] = wireIn[147];    
  assign wireOut[167] = wireIn[211];    
  assign wireOut[168] = wireIn[148];    
  assign wireOut[169] = wireIn[212];    
  assign wireOut[170] = wireIn[149];    
  assign wireOut[171] = wireIn[213];    
  assign wireOut[172] = wireIn[150];    
  assign wireOut[173] = wireIn[214];    
  assign wireOut[174] = wireIn[151];    
  assign wireOut[175] = wireIn[215];    
  assign wireOut[176] = wireIn[152];    
  assign wireOut[177] = wireIn[216];    
  assign wireOut[178] = wireIn[153];    
  assign wireOut[179] = wireIn[217];    
  assign wireOut[180] = wireIn[154];    
  assign wireOut[181] = wireIn[218];    
  assign wireOut[182] = wireIn[155];    
  assign wireOut[183] = wireIn[219];    
  assign wireOut[184] = wireIn[156];    
  assign wireOut[185] = wireIn[220];    
  assign wireOut[186] = wireIn[157];    
  assign wireOut[187] = wireIn[221];    
  assign wireOut[188] = wireIn[158];    
  assign wireOut[189] = wireIn[222];    
  assign wireOut[190] = wireIn[159];    
  assign wireOut[191] = wireIn[223];    
  assign wireOut[192] = wireIn[160];    
  assign wireOut[193] = wireIn[224];    
  assign wireOut[194] = wireIn[161];    
  assign wireOut[195] = wireIn[225];    
  assign wireOut[196] = wireIn[162];    
  assign wireOut[197] = wireIn[226];    
  assign wireOut[198] = wireIn[163];    
  assign wireOut[199] = wireIn[227];    
  assign wireOut[200] = wireIn[164];    
  assign wireOut[201] = wireIn[228];    
  assign wireOut[202] = wireIn[165];    
  assign wireOut[203] = wireIn[229];    
  assign wireOut[204] = wireIn[166];    
  assign wireOut[205] = wireIn[230];    
  assign wireOut[206] = wireIn[167];    
  assign wireOut[207] = wireIn[231];    
  assign wireOut[208] = wireIn[168];    
  assign wireOut[209] = wireIn[232];    
  assign wireOut[210] = wireIn[169];    
  assign wireOut[211] = wireIn[233];    
  assign wireOut[212] = wireIn[170];    
  assign wireOut[213] = wireIn[234];    
  assign wireOut[214] = wireIn[171];    
  assign wireOut[215] = wireIn[235];    
  assign wireOut[216] = wireIn[172];    
  assign wireOut[217] = wireIn[236];    
  assign wireOut[218] = wireIn[173];    
  assign wireOut[219] = wireIn[237];    
  assign wireOut[220] = wireIn[174];    
  assign wireOut[221] = wireIn[238];    
  assign wireOut[222] = wireIn[175];    
  assign wireOut[223] = wireIn[239];    
  assign wireOut[224] = wireIn[176];    
  assign wireOut[225] = wireIn[240];    
  assign wireOut[226] = wireIn[177];    
  assign wireOut[227] = wireIn[241];    
  assign wireOut[228] = wireIn[178];    
  assign wireOut[229] = wireIn[242];    
  assign wireOut[230] = wireIn[179];    
  assign wireOut[231] = wireIn[243];    
  assign wireOut[232] = wireIn[180];    
  assign wireOut[233] = wireIn[244];    
  assign wireOut[234] = wireIn[181];    
  assign wireOut[235] = wireIn[245];    
  assign wireOut[236] = wireIn[182];    
  assign wireOut[237] = wireIn[246];    
  assign wireOut[238] = wireIn[183];    
  assign wireOut[239] = wireIn[247];    
  assign wireOut[240] = wireIn[184];    
  assign wireOut[241] = wireIn[248];    
  assign wireOut[242] = wireIn[185];    
  assign wireOut[243] = wireIn[249];    
  assign wireOut[244] = wireIn[186];    
  assign wireOut[245] = wireIn[250];    
  assign wireOut[246] = wireIn[187];    
  assign wireOut[247] = wireIn[251];    
  assign wireOut[248] = wireIn[188];    
  assign wireOut[249] = wireIn[252];    
  assign wireOut[250] = wireIn[189];    
  assign wireOut[251] = wireIn[253];    
  assign wireOut[252] = wireIn[190];    
  assign wireOut[253] = wireIn[254];    
  assign wireOut[254] = wireIn[191];    
  assign wireOut[255] = wireIn[255];    
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module switches_stage_st2_0_R(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
ctrl,                            
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;                   
  input [128-1:0] ctrl;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  switch_2_2 switch_inst_0(.inData_0(wireIn[0]), .inData_1(wireIn[1]), .outData_0(wireOut[0]), .outData_1(wireOut[1]), .ctrl(ctrl[0]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_1(.inData_0(wireIn[2]), .inData_1(wireIn[3]), .outData_0(wireOut[2]), .outData_1(wireOut[3]), .ctrl(ctrl[1]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_2(.inData_0(wireIn[4]), .inData_1(wireIn[5]), .outData_0(wireOut[4]), .outData_1(wireOut[5]), .ctrl(ctrl[2]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_3(.inData_0(wireIn[6]), .inData_1(wireIn[7]), .outData_0(wireOut[6]), .outData_1(wireOut[7]), .ctrl(ctrl[3]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_4(.inData_0(wireIn[8]), .inData_1(wireIn[9]), .outData_0(wireOut[8]), .outData_1(wireOut[9]), .ctrl(ctrl[4]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_5(.inData_0(wireIn[10]), .inData_1(wireIn[11]), .outData_0(wireOut[10]), .outData_1(wireOut[11]), .ctrl(ctrl[5]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_6(.inData_0(wireIn[12]), .inData_1(wireIn[13]), .outData_0(wireOut[12]), .outData_1(wireOut[13]), .ctrl(ctrl[6]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_7(.inData_0(wireIn[14]), .inData_1(wireIn[15]), .outData_0(wireOut[14]), .outData_1(wireOut[15]), .ctrl(ctrl[7]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_8(.inData_0(wireIn[16]), .inData_1(wireIn[17]), .outData_0(wireOut[16]), .outData_1(wireOut[17]), .ctrl(ctrl[8]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_9(.inData_0(wireIn[18]), .inData_1(wireIn[19]), .outData_0(wireOut[18]), .outData_1(wireOut[19]), .ctrl(ctrl[9]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_10(.inData_0(wireIn[20]), .inData_1(wireIn[21]), .outData_0(wireOut[20]), .outData_1(wireOut[21]), .ctrl(ctrl[10]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_11(.inData_0(wireIn[22]), .inData_1(wireIn[23]), .outData_0(wireOut[22]), .outData_1(wireOut[23]), .ctrl(ctrl[11]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_12(.inData_0(wireIn[24]), .inData_1(wireIn[25]), .outData_0(wireOut[24]), .outData_1(wireOut[25]), .ctrl(ctrl[12]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_13(.inData_0(wireIn[26]), .inData_1(wireIn[27]), .outData_0(wireOut[26]), .outData_1(wireOut[27]), .ctrl(ctrl[13]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_14(.inData_0(wireIn[28]), .inData_1(wireIn[29]), .outData_0(wireOut[28]), .outData_1(wireOut[29]), .ctrl(ctrl[14]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_15(.inData_0(wireIn[30]), .inData_1(wireIn[31]), .outData_0(wireOut[30]), .outData_1(wireOut[31]), .ctrl(ctrl[15]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_16(.inData_0(wireIn[32]), .inData_1(wireIn[33]), .outData_0(wireOut[32]), .outData_1(wireOut[33]), .ctrl(ctrl[16]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_17(.inData_0(wireIn[34]), .inData_1(wireIn[35]), .outData_0(wireOut[34]), .outData_1(wireOut[35]), .ctrl(ctrl[17]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_18(.inData_0(wireIn[36]), .inData_1(wireIn[37]), .outData_0(wireOut[36]), .outData_1(wireOut[37]), .ctrl(ctrl[18]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_19(.inData_0(wireIn[38]), .inData_1(wireIn[39]), .outData_0(wireOut[38]), .outData_1(wireOut[39]), .ctrl(ctrl[19]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_20(.inData_0(wireIn[40]), .inData_1(wireIn[41]), .outData_0(wireOut[40]), .outData_1(wireOut[41]), .ctrl(ctrl[20]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_21(.inData_0(wireIn[42]), .inData_1(wireIn[43]), .outData_0(wireOut[42]), .outData_1(wireOut[43]), .ctrl(ctrl[21]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_22(.inData_0(wireIn[44]), .inData_1(wireIn[45]), .outData_0(wireOut[44]), .outData_1(wireOut[45]), .ctrl(ctrl[22]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_23(.inData_0(wireIn[46]), .inData_1(wireIn[47]), .outData_0(wireOut[46]), .outData_1(wireOut[47]), .ctrl(ctrl[23]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_24(.inData_0(wireIn[48]), .inData_1(wireIn[49]), .outData_0(wireOut[48]), .outData_1(wireOut[49]), .ctrl(ctrl[24]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_25(.inData_0(wireIn[50]), .inData_1(wireIn[51]), .outData_0(wireOut[50]), .outData_1(wireOut[51]), .ctrl(ctrl[25]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_26(.inData_0(wireIn[52]), .inData_1(wireIn[53]), .outData_0(wireOut[52]), .outData_1(wireOut[53]), .ctrl(ctrl[26]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_27(.inData_0(wireIn[54]), .inData_1(wireIn[55]), .outData_0(wireOut[54]), .outData_1(wireOut[55]), .ctrl(ctrl[27]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_28(.inData_0(wireIn[56]), .inData_1(wireIn[57]), .outData_0(wireOut[56]), .outData_1(wireOut[57]), .ctrl(ctrl[28]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_29(.inData_0(wireIn[58]), .inData_1(wireIn[59]), .outData_0(wireOut[58]), .outData_1(wireOut[59]), .ctrl(ctrl[29]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_30(.inData_0(wireIn[60]), .inData_1(wireIn[61]), .outData_0(wireOut[60]), .outData_1(wireOut[61]), .ctrl(ctrl[30]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_31(.inData_0(wireIn[62]), .inData_1(wireIn[63]), .outData_0(wireOut[62]), .outData_1(wireOut[63]), .ctrl(ctrl[31]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_32(.inData_0(wireIn[64]), .inData_1(wireIn[65]), .outData_0(wireOut[64]), .outData_1(wireOut[65]), .ctrl(ctrl[32]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_33(.inData_0(wireIn[66]), .inData_1(wireIn[67]), .outData_0(wireOut[66]), .outData_1(wireOut[67]), .ctrl(ctrl[33]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_34(.inData_0(wireIn[68]), .inData_1(wireIn[69]), .outData_0(wireOut[68]), .outData_1(wireOut[69]), .ctrl(ctrl[34]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_35(.inData_0(wireIn[70]), .inData_1(wireIn[71]), .outData_0(wireOut[70]), .outData_1(wireOut[71]), .ctrl(ctrl[35]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_36(.inData_0(wireIn[72]), .inData_1(wireIn[73]), .outData_0(wireOut[72]), .outData_1(wireOut[73]), .ctrl(ctrl[36]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_37(.inData_0(wireIn[74]), .inData_1(wireIn[75]), .outData_0(wireOut[74]), .outData_1(wireOut[75]), .ctrl(ctrl[37]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_38(.inData_0(wireIn[76]), .inData_1(wireIn[77]), .outData_0(wireOut[76]), .outData_1(wireOut[77]), .ctrl(ctrl[38]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_39(.inData_0(wireIn[78]), .inData_1(wireIn[79]), .outData_0(wireOut[78]), .outData_1(wireOut[79]), .ctrl(ctrl[39]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_40(.inData_0(wireIn[80]), .inData_1(wireIn[81]), .outData_0(wireOut[80]), .outData_1(wireOut[81]), .ctrl(ctrl[40]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_41(.inData_0(wireIn[82]), .inData_1(wireIn[83]), .outData_0(wireOut[82]), .outData_1(wireOut[83]), .ctrl(ctrl[41]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_42(.inData_0(wireIn[84]), .inData_1(wireIn[85]), .outData_0(wireOut[84]), .outData_1(wireOut[85]), .ctrl(ctrl[42]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_43(.inData_0(wireIn[86]), .inData_1(wireIn[87]), .outData_0(wireOut[86]), .outData_1(wireOut[87]), .ctrl(ctrl[43]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_44(.inData_0(wireIn[88]), .inData_1(wireIn[89]), .outData_0(wireOut[88]), .outData_1(wireOut[89]), .ctrl(ctrl[44]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_45(.inData_0(wireIn[90]), .inData_1(wireIn[91]), .outData_0(wireOut[90]), .outData_1(wireOut[91]), .ctrl(ctrl[45]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_46(.inData_0(wireIn[92]), .inData_1(wireIn[93]), .outData_0(wireOut[92]), .outData_1(wireOut[93]), .ctrl(ctrl[46]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_47(.inData_0(wireIn[94]), .inData_1(wireIn[95]), .outData_0(wireOut[94]), .outData_1(wireOut[95]), .ctrl(ctrl[47]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_48(.inData_0(wireIn[96]), .inData_1(wireIn[97]), .outData_0(wireOut[96]), .outData_1(wireOut[97]), .ctrl(ctrl[48]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_49(.inData_0(wireIn[98]), .inData_1(wireIn[99]), .outData_0(wireOut[98]), .outData_1(wireOut[99]), .ctrl(ctrl[49]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_50(.inData_0(wireIn[100]), .inData_1(wireIn[101]), .outData_0(wireOut[100]), .outData_1(wireOut[101]), .ctrl(ctrl[50]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_51(.inData_0(wireIn[102]), .inData_1(wireIn[103]), .outData_0(wireOut[102]), .outData_1(wireOut[103]), .ctrl(ctrl[51]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_52(.inData_0(wireIn[104]), .inData_1(wireIn[105]), .outData_0(wireOut[104]), .outData_1(wireOut[105]), .ctrl(ctrl[52]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_53(.inData_0(wireIn[106]), .inData_1(wireIn[107]), .outData_0(wireOut[106]), .outData_1(wireOut[107]), .ctrl(ctrl[53]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_54(.inData_0(wireIn[108]), .inData_1(wireIn[109]), .outData_0(wireOut[108]), .outData_1(wireOut[109]), .ctrl(ctrl[54]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_55(.inData_0(wireIn[110]), .inData_1(wireIn[111]), .outData_0(wireOut[110]), .outData_1(wireOut[111]), .ctrl(ctrl[55]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_56(.inData_0(wireIn[112]), .inData_1(wireIn[113]), .outData_0(wireOut[112]), .outData_1(wireOut[113]), .ctrl(ctrl[56]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_57(.inData_0(wireIn[114]), .inData_1(wireIn[115]), .outData_0(wireOut[114]), .outData_1(wireOut[115]), .ctrl(ctrl[57]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_58(.inData_0(wireIn[116]), .inData_1(wireIn[117]), .outData_0(wireOut[116]), .outData_1(wireOut[117]), .ctrl(ctrl[58]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_59(.inData_0(wireIn[118]), .inData_1(wireIn[119]), .outData_0(wireOut[118]), .outData_1(wireOut[119]), .ctrl(ctrl[59]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_60(.inData_0(wireIn[120]), .inData_1(wireIn[121]), .outData_0(wireOut[120]), .outData_1(wireOut[121]), .ctrl(ctrl[60]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_61(.inData_0(wireIn[122]), .inData_1(wireIn[123]), .outData_0(wireOut[122]), .outData_1(wireOut[123]), .ctrl(ctrl[61]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_62(.inData_0(wireIn[124]), .inData_1(wireIn[125]), .outData_0(wireOut[124]), .outData_1(wireOut[125]), .ctrl(ctrl[62]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_63(.inData_0(wireIn[126]), .inData_1(wireIn[127]), .outData_0(wireOut[126]), .outData_1(wireOut[127]), .ctrl(ctrl[63]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_64(.inData_0(wireIn[128]), .inData_1(wireIn[129]), .outData_0(wireOut[128]), .outData_1(wireOut[129]), .ctrl(ctrl[64]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_65(.inData_0(wireIn[130]), .inData_1(wireIn[131]), .outData_0(wireOut[130]), .outData_1(wireOut[131]), .ctrl(ctrl[65]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_66(.inData_0(wireIn[132]), .inData_1(wireIn[133]), .outData_0(wireOut[132]), .outData_1(wireOut[133]), .ctrl(ctrl[66]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_67(.inData_0(wireIn[134]), .inData_1(wireIn[135]), .outData_0(wireOut[134]), .outData_1(wireOut[135]), .ctrl(ctrl[67]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_68(.inData_0(wireIn[136]), .inData_1(wireIn[137]), .outData_0(wireOut[136]), .outData_1(wireOut[137]), .ctrl(ctrl[68]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_69(.inData_0(wireIn[138]), .inData_1(wireIn[139]), .outData_0(wireOut[138]), .outData_1(wireOut[139]), .ctrl(ctrl[69]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_70(.inData_0(wireIn[140]), .inData_1(wireIn[141]), .outData_0(wireOut[140]), .outData_1(wireOut[141]), .ctrl(ctrl[70]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_71(.inData_0(wireIn[142]), .inData_1(wireIn[143]), .outData_0(wireOut[142]), .outData_1(wireOut[143]), .ctrl(ctrl[71]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_72(.inData_0(wireIn[144]), .inData_1(wireIn[145]), .outData_0(wireOut[144]), .outData_1(wireOut[145]), .ctrl(ctrl[72]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_73(.inData_0(wireIn[146]), .inData_1(wireIn[147]), .outData_0(wireOut[146]), .outData_1(wireOut[147]), .ctrl(ctrl[73]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_74(.inData_0(wireIn[148]), .inData_1(wireIn[149]), .outData_0(wireOut[148]), .outData_1(wireOut[149]), .ctrl(ctrl[74]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_75(.inData_0(wireIn[150]), .inData_1(wireIn[151]), .outData_0(wireOut[150]), .outData_1(wireOut[151]), .ctrl(ctrl[75]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_76(.inData_0(wireIn[152]), .inData_1(wireIn[153]), .outData_0(wireOut[152]), .outData_1(wireOut[153]), .ctrl(ctrl[76]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_77(.inData_0(wireIn[154]), .inData_1(wireIn[155]), .outData_0(wireOut[154]), .outData_1(wireOut[155]), .ctrl(ctrl[77]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_78(.inData_0(wireIn[156]), .inData_1(wireIn[157]), .outData_0(wireOut[156]), .outData_1(wireOut[157]), .ctrl(ctrl[78]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_79(.inData_0(wireIn[158]), .inData_1(wireIn[159]), .outData_0(wireOut[158]), .outData_1(wireOut[159]), .ctrl(ctrl[79]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_80(.inData_0(wireIn[160]), .inData_1(wireIn[161]), .outData_0(wireOut[160]), .outData_1(wireOut[161]), .ctrl(ctrl[80]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_81(.inData_0(wireIn[162]), .inData_1(wireIn[163]), .outData_0(wireOut[162]), .outData_1(wireOut[163]), .ctrl(ctrl[81]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_82(.inData_0(wireIn[164]), .inData_1(wireIn[165]), .outData_0(wireOut[164]), .outData_1(wireOut[165]), .ctrl(ctrl[82]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_83(.inData_0(wireIn[166]), .inData_1(wireIn[167]), .outData_0(wireOut[166]), .outData_1(wireOut[167]), .ctrl(ctrl[83]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_84(.inData_0(wireIn[168]), .inData_1(wireIn[169]), .outData_0(wireOut[168]), .outData_1(wireOut[169]), .ctrl(ctrl[84]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_85(.inData_0(wireIn[170]), .inData_1(wireIn[171]), .outData_0(wireOut[170]), .outData_1(wireOut[171]), .ctrl(ctrl[85]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_86(.inData_0(wireIn[172]), .inData_1(wireIn[173]), .outData_0(wireOut[172]), .outData_1(wireOut[173]), .ctrl(ctrl[86]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_87(.inData_0(wireIn[174]), .inData_1(wireIn[175]), .outData_0(wireOut[174]), .outData_1(wireOut[175]), .ctrl(ctrl[87]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_88(.inData_0(wireIn[176]), .inData_1(wireIn[177]), .outData_0(wireOut[176]), .outData_1(wireOut[177]), .ctrl(ctrl[88]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_89(.inData_0(wireIn[178]), .inData_1(wireIn[179]), .outData_0(wireOut[178]), .outData_1(wireOut[179]), .ctrl(ctrl[89]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_90(.inData_0(wireIn[180]), .inData_1(wireIn[181]), .outData_0(wireOut[180]), .outData_1(wireOut[181]), .ctrl(ctrl[90]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_91(.inData_0(wireIn[182]), .inData_1(wireIn[183]), .outData_0(wireOut[182]), .outData_1(wireOut[183]), .ctrl(ctrl[91]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_92(.inData_0(wireIn[184]), .inData_1(wireIn[185]), .outData_0(wireOut[184]), .outData_1(wireOut[185]), .ctrl(ctrl[92]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_93(.inData_0(wireIn[186]), .inData_1(wireIn[187]), .outData_0(wireOut[186]), .outData_1(wireOut[187]), .ctrl(ctrl[93]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_94(.inData_0(wireIn[188]), .inData_1(wireIn[189]), .outData_0(wireOut[188]), .outData_1(wireOut[189]), .ctrl(ctrl[94]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_95(.inData_0(wireIn[190]), .inData_1(wireIn[191]), .outData_0(wireOut[190]), .outData_1(wireOut[191]), .ctrl(ctrl[95]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_96(.inData_0(wireIn[192]), .inData_1(wireIn[193]), .outData_0(wireOut[192]), .outData_1(wireOut[193]), .ctrl(ctrl[96]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_97(.inData_0(wireIn[194]), .inData_1(wireIn[195]), .outData_0(wireOut[194]), .outData_1(wireOut[195]), .ctrl(ctrl[97]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_98(.inData_0(wireIn[196]), .inData_1(wireIn[197]), .outData_0(wireOut[196]), .outData_1(wireOut[197]), .ctrl(ctrl[98]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_99(.inData_0(wireIn[198]), .inData_1(wireIn[199]), .outData_0(wireOut[198]), .outData_1(wireOut[199]), .ctrl(ctrl[99]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_100(.inData_0(wireIn[200]), .inData_1(wireIn[201]), .outData_0(wireOut[200]), .outData_1(wireOut[201]), .ctrl(ctrl[100]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_101(.inData_0(wireIn[202]), .inData_1(wireIn[203]), .outData_0(wireOut[202]), .outData_1(wireOut[203]), .ctrl(ctrl[101]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_102(.inData_0(wireIn[204]), .inData_1(wireIn[205]), .outData_0(wireOut[204]), .outData_1(wireOut[205]), .ctrl(ctrl[102]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_103(.inData_0(wireIn[206]), .inData_1(wireIn[207]), .outData_0(wireOut[206]), .outData_1(wireOut[207]), .ctrl(ctrl[103]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_104(.inData_0(wireIn[208]), .inData_1(wireIn[209]), .outData_0(wireOut[208]), .outData_1(wireOut[209]), .ctrl(ctrl[104]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_105(.inData_0(wireIn[210]), .inData_1(wireIn[211]), .outData_0(wireOut[210]), .outData_1(wireOut[211]), .ctrl(ctrl[105]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_106(.inData_0(wireIn[212]), .inData_1(wireIn[213]), .outData_0(wireOut[212]), .outData_1(wireOut[213]), .ctrl(ctrl[106]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_107(.inData_0(wireIn[214]), .inData_1(wireIn[215]), .outData_0(wireOut[214]), .outData_1(wireOut[215]), .ctrl(ctrl[107]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_108(.inData_0(wireIn[216]), .inData_1(wireIn[217]), .outData_0(wireOut[216]), .outData_1(wireOut[217]), .ctrl(ctrl[108]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_109(.inData_0(wireIn[218]), .inData_1(wireIn[219]), .outData_0(wireOut[218]), .outData_1(wireOut[219]), .ctrl(ctrl[109]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_110(.inData_0(wireIn[220]), .inData_1(wireIn[221]), .outData_0(wireOut[220]), .outData_1(wireOut[221]), .ctrl(ctrl[110]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_111(.inData_0(wireIn[222]), .inData_1(wireIn[223]), .outData_0(wireOut[222]), .outData_1(wireOut[223]), .ctrl(ctrl[111]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_112(.inData_0(wireIn[224]), .inData_1(wireIn[225]), .outData_0(wireOut[224]), .outData_1(wireOut[225]), .ctrl(ctrl[112]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_113(.inData_0(wireIn[226]), .inData_1(wireIn[227]), .outData_0(wireOut[226]), .outData_1(wireOut[227]), .ctrl(ctrl[113]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_114(.inData_0(wireIn[228]), .inData_1(wireIn[229]), .outData_0(wireOut[228]), .outData_1(wireOut[229]), .ctrl(ctrl[114]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_115(.inData_0(wireIn[230]), .inData_1(wireIn[231]), .outData_0(wireOut[230]), .outData_1(wireOut[231]), .ctrl(ctrl[115]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_116(.inData_0(wireIn[232]), .inData_1(wireIn[233]), .outData_0(wireOut[232]), .outData_1(wireOut[233]), .ctrl(ctrl[116]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_117(.inData_0(wireIn[234]), .inData_1(wireIn[235]), .outData_0(wireOut[234]), .outData_1(wireOut[235]), .ctrl(ctrl[117]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_118(.inData_0(wireIn[236]), .inData_1(wireIn[237]), .outData_0(wireOut[236]), .outData_1(wireOut[237]), .ctrl(ctrl[118]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_119(.inData_0(wireIn[238]), .inData_1(wireIn[239]), .outData_0(wireOut[238]), .outData_1(wireOut[239]), .ctrl(ctrl[119]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_120(.inData_0(wireIn[240]), .inData_1(wireIn[241]), .outData_0(wireOut[240]), .outData_1(wireOut[241]), .ctrl(ctrl[120]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_121(.inData_0(wireIn[242]), .inData_1(wireIn[243]), .outData_0(wireOut[242]), .outData_1(wireOut[243]), .ctrl(ctrl[121]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_122(.inData_0(wireIn[244]), .inData_1(wireIn[245]), .outData_0(wireOut[244]), .outData_1(wireOut[245]), .ctrl(ctrl[122]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_123(.inData_0(wireIn[246]), .inData_1(wireIn[247]), .outData_0(wireOut[246]), .outData_1(wireOut[247]), .ctrl(ctrl[123]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_124(.inData_0(wireIn[248]), .inData_1(wireIn[249]), .outData_0(wireOut[248]), .outData_1(wireOut[249]), .ctrl(ctrl[124]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_125(.inData_0(wireIn[250]), .inData_1(wireIn[251]), .outData_0(wireOut[250]), .outData_1(wireOut[251]), .ctrl(ctrl[125]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_126(.inData_0(wireIn[252]), .inData_1(wireIn[253]), .outData_0(wireOut[252]), .outData_1(wireOut[253]), .ctrl(ctrl[126]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_127(.inData_0(wireIn[254]), .inData_1(wireIn[255]), .outData_0(wireOut[254]), .outData_1(wireOut[255]), .ctrl(ctrl[127]), .clk(clk), .rst(rst));
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module wireCon_dp256_st2_R(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  assign wireOut[0] = wireIn[0];    
  assign wireOut[1] = wireIn[32];    
  assign wireOut[2] = wireIn[1];    
  assign wireOut[3] = wireIn[33];    
  assign wireOut[4] = wireIn[2];    
  assign wireOut[5] = wireIn[34];    
  assign wireOut[6] = wireIn[3];    
  assign wireOut[7] = wireIn[35];    
  assign wireOut[8] = wireIn[4];    
  assign wireOut[9] = wireIn[36];    
  assign wireOut[10] = wireIn[5];    
  assign wireOut[11] = wireIn[37];    
  assign wireOut[12] = wireIn[6];    
  assign wireOut[13] = wireIn[38];    
  assign wireOut[14] = wireIn[7];    
  assign wireOut[15] = wireIn[39];    
  assign wireOut[16] = wireIn[8];    
  assign wireOut[17] = wireIn[40];    
  assign wireOut[18] = wireIn[9];    
  assign wireOut[19] = wireIn[41];    
  assign wireOut[20] = wireIn[10];    
  assign wireOut[21] = wireIn[42];    
  assign wireOut[22] = wireIn[11];    
  assign wireOut[23] = wireIn[43];    
  assign wireOut[24] = wireIn[12];    
  assign wireOut[25] = wireIn[44];    
  assign wireOut[26] = wireIn[13];    
  assign wireOut[27] = wireIn[45];    
  assign wireOut[28] = wireIn[14];    
  assign wireOut[29] = wireIn[46];    
  assign wireOut[30] = wireIn[15];    
  assign wireOut[31] = wireIn[47];    
  assign wireOut[32] = wireIn[16];    
  assign wireOut[33] = wireIn[48];    
  assign wireOut[34] = wireIn[17];    
  assign wireOut[35] = wireIn[49];    
  assign wireOut[36] = wireIn[18];    
  assign wireOut[37] = wireIn[50];    
  assign wireOut[38] = wireIn[19];    
  assign wireOut[39] = wireIn[51];    
  assign wireOut[40] = wireIn[20];    
  assign wireOut[41] = wireIn[52];    
  assign wireOut[42] = wireIn[21];    
  assign wireOut[43] = wireIn[53];    
  assign wireOut[44] = wireIn[22];    
  assign wireOut[45] = wireIn[54];    
  assign wireOut[46] = wireIn[23];    
  assign wireOut[47] = wireIn[55];    
  assign wireOut[48] = wireIn[24];    
  assign wireOut[49] = wireIn[56];    
  assign wireOut[50] = wireIn[25];    
  assign wireOut[51] = wireIn[57];    
  assign wireOut[52] = wireIn[26];    
  assign wireOut[53] = wireIn[58];    
  assign wireOut[54] = wireIn[27];    
  assign wireOut[55] = wireIn[59];    
  assign wireOut[56] = wireIn[28];    
  assign wireOut[57] = wireIn[60];    
  assign wireOut[58] = wireIn[29];    
  assign wireOut[59] = wireIn[61];    
  assign wireOut[60] = wireIn[30];    
  assign wireOut[61] = wireIn[62];    
  assign wireOut[62] = wireIn[31];    
  assign wireOut[63] = wireIn[63];    
  assign wireOut[64] = wireIn[64];    
  assign wireOut[65] = wireIn[96];    
  assign wireOut[66] = wireIn[65];    
  assign wireOut[67] = wireIn[97];    
  assign wireOut[68] = wireIn[66];    
  assign wireOut[69] = wireIn[98];    
  assign wireOut[70] = wireIn[67];    
  assign wireOut[71] = wireIn[99];    
  assign wireOut[72] = wireIn[68];    
  assign wireOut[73] = wireIn[100];    
  assign wireOut[74] = wireIn[69];    
  assign wireOut[75] = wireIn[101];    
  assign wireOut[76] = wireIn[70];    
  assign wireOut[77] = wireIn[102];    
  assign wireOut[78] = wireIn[71];    
  assign wireOut[79] = wireIn[103];    
  assign wireOut[80] = wireIn[72];    
  assign wireOut[81] = wireIn[104];    
  assign wireOut[82] = wireIn[73];    
  assign wireOut[83] = wireIn[105];    
  assign wireOut[84] = wireIn[74];    
  assign wireOut[85] = wireIn[106];    
  assign wireOut[86] = wireIn[75];    
  assign wireOut[87] = wireIn[107];    
  assign wireOut[88] = wireIn[76];    
  assign wireOut[89] = wireIn[108];    
  assign wireOut[90] = wireIn[77];    
  assign wireOut[91] = wireIn[109];    
  assign wireOut[92] = wireIn[78];    
  assign wireOut[93] = wireIn[110];    
  assign wireOut[94] = wireIn[79];    
  assign wireOut[95] = wireIn[111];    
  assign wireOut[96] = wireIn[80];    
  assign wireOut[97] = wireIn[112];    
  assign wireOut[98] = wireIn[81];    
  assign wireOut[99] = wireIn[113];    
  assign wireOut[100] = wireIn[82];    
  assign wireOut[101] = wireIn[114];    
  assign wireOut[102] = wireIn[83];    
  assign wireOut[103] = wireIn[115];    
  assign wireOut[104] = wireIn[84];    
  assign wireOut[105] = wireIn[116];    
  assign wireOut[106] = wireIn[85];    
  assign wireOut[107] = wireIn[117];    
  assign wireOut[108] = wireIn[86];    
  assign wireOut[109] = wireIn[118];    
  assign wireOut[110] = wireIn[87];    
  assign wireOut[111] = wireIn[119];    
  assign wireOut[112] = wireIn[88];    
  assign wireOut[113] = wireIn[120];    
  assign wireOut[114] = wireIn[89];    
  assign wireOut[115] = wireIn[121];    
  assign wireOut[116] = wireIn[90];    
  assign wireOut[117] = wireIn[122];    
  assign wireOut[118] = wireIn[91];    
  assign wireOut[119] = wireIn[123];    
  assign wireOut[120] = wireIn[92];    
  assign wireOut[121] = wireIn[124];    
  assign wireOut[122] = wireIn[93];    
  assign wireOut[123] = wireIn[125];    
  assign wireOut[124] = wireIn[94];    
  assign wireOut[125] = wireIn[126];    
  assign wireOut[126] = wireIn[95];    
  assign wireOut[127] = wireIn[127];    
  assign wireOut[128] = wireIn[128];    
  assign wireOut[129] = wireIn[160];    
  assign wireOut[130] = wireIn[129];    
  assign wireOut[131] = wireIn[161];    
  assign wireOut[132] = wireIn[130];    
  assign wireOut[133] = wireIn[162];    
  assign wireOut[134] = wireIn[131];    
  assign wireOut[135] = wireIn[163];    
  assign wireOut[136] = wireIn[132];    
  assign wireOut[137] = wireIn[164];    
  assign wireOut[138] = wireIn[133];    
  assign wireOut[139] = wireIn[165];    
  assign wireOut[140] = wireIn[134];    
  assign wireOut[141] = wireIn[166];    
  assign wireOut[142] = wireIn[135];    
  assign wireOut[143] = wireIn[167];    
  assign wireOut[144] = wireIn[136];    
  assign wireOut[145] = wireIn[168];    
  assign wireOut[146] = wireIn[137];    
  assign wireOut[147] = wireIn[169];    
  assign wireOut[148] = wireIn[138];    
  assign wireOut[149] = wireIn[170];    
  assign wireOut[150] = wireIn[139];    
  assign wireOut[151] = wireIn[171];    
  assign wireOut[152] = wireIn[140];    
  assign wireOut[153] = wireIn[172];    
  assign wireOut[154] = wireIn[141];    
  assign wireOut[155] = wireIn[173];    
  assign wireOut[156] = wireIn[142];    
  assign wireOut[157] = wireIn[174];    
  assign wireOut[158] = wireIn[143];    
  assign wireOut[159] = wireIn[175];    
  assign wireOut[160] = wireIn[144];    
  assign wireOut[161] = wireIn[176];    
  assign wireOut[162] = wireIn[145];    
  assign wireOut[163] = wireIn[177];    
  assign wireOut[164] = wireIn[146];    
  assign wireOut[165] = wireIn[178];    
  assign wireOut[166] = wireIn[147];    
  assign wireOut[167] = wireIn[179];    
  assign wireOut[168] = wireIn[148];    
  assign wireOut[169] = wireIn[180];    
  assign wireOut[170] = wireIn[149];    
  assign wireOut[171] = wireIn[181];    
  assign wireOut[172] = wireIn[150];    
  assign wireOut[173] = wireIn[182];    
  assign wireOut[174] = wireIn[151];    
  assign wireOut[175] = wireIn[183];    
  assign wireOut[176] = wireIn[152];    
  assign wireOut[177] = wireIn[184];    
  assign wireOut[178] = wireIn[153];    
  assign wireOut[179] = wireIn[185];    
  assign wireOut[180] = wireIn[154];    
  assign wireOut[181] = wireIn[186];    
  assign wireOut[182] = wireIn[155];    
  assign wireOut[183] = wireIn[187];    
  assign wireOut[184] = wireIn[156];    
  assign wireOut[185] = wireIn[188];    
  assign wireOut[186] = wireIn[157];    
  assign wireOut[187] = wireIn[189];    
  assign wireOut[188] = wireIn[158];    
  assign wireOut[189] = wireIn[190];    
  assign wireOut[190] = wireIn[159];    
  assign wireOut[191] = wireIn[191];    
  assign wireOut[192] = wireIn[192];    
  assign wireOut[193] = wireIn[224];    
  assign wireOut[194] = wireIn[193];    
  assign wireOut[195] = wireIn[225];    
  assign wireOut[196] = wireIn[194];    
  assign wireOut[197] = wireIn[226];    
  assign wireOut[198] = wireIn[195];    
  assign wireOut[199] = wireIn[227];    
  assign wireOut[200] = wireIn[196];    
  assign wireOut[201] = wireIn[228];    
  assign wireOut[202] = wireIn[197];    
  assign wireOut[203] = wireIn[229];    
  assign wireOut[204] = wireIn[198];    
  assign wireOut[205] = wireIn[230];    
  assign wireOut[206] = wireIn[199];    
  assign wireOut[207] = wireIn[231];    
  assign wireOut[208] = wireIn[200];    
  assign wireOut[209] = wireIn[232];    
  assign wireOut[210] = wireIn[201];    
  assign wireOut[211] = wireIn[233];    
  assign wireOut[212] = wireIn[202];    
  assign wireOut[213] = wireIn[234];    
  assign wireOut[214] = wireIn[203];    
  assign wireOut[215] = wireIn[235];    
  assign wireOut[216] = wireIn[204];    
  assign wireOut[217] = wireIn[236];    
  assign wireOut[218] = wireIn[205];    
  assign wireOut[219] = wireIn[237];    
  assign wireOut[220] = wireIn[206];    
  assign wireOut[221] = wireIn[238];    
  assign wireOut[222] = wireIn[207];    
  assign wireOut[223] = wireIn[239];    
  assign wireOut[224] = wireIn[208];    
  assign wireOut[225] = wireIn[240];    
  assign wireOut[226] = wireIn[209];    
  assign wireOut[227] = wireIn[241];    
  assign wireOut[228] = wireIn[210];    
  assign wireOut[229] = wireIn[242];    
  assign wireOut[230] = wireIn[211];    
  assign wireOut[231] = wireIn[243];    
  assign wireOut[232] = wireIn[212];    
  assign wireOut[233] = wireIn[244];    
  assign wireOut[234] = wireIn[213];    
  assign wireOut[235] = wireIn[245];    
  assign wireOut[236] = wireIn[214];    
  assign wireOut[237] = wireIn[246];    
  assign wireOut[238] = wireIn[215];    
  assign wireOut[239] = wireIn[247];    
  assign wireOut[240] = wireIn[216];    
  assign wireOut[241] = wireIn[248];    
  assign wireOut[242] = wireIn[217];    
  assign wireOut[243] = wireIn[249];    
  assign wireOut[244] = wireIn[218];    
  assign wireOut[245] = wireIn[250];    
  assign wireOut[246] = wireIn[219];    
  assign wireOut[247] = wireIn[251];    
  assign wireOut[248] = wireIn[220];    
  assign wireOut[249] = wireIn[252];    
  assign wireOut[250] = wireIn[221];    
  assign wireOut[251] = wireIn[253];    
  assign wireOut[252] = wireIn[222];    
  assign wireOut[253] = wireIn[254];    
  assign wireOut[254] = wireIn[223];    
  assign wireOut[255] = wireIn[255];    
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module switches_stage_st3_0_R(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
ctrl,                            
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;                   
  input [128-1:0] ctrl;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  switch_2_2 switch_inst_0(.inData_0(wireIn[0]), .inData_1(wireIn[1]), .outData_0(wireOut[0]), .outData_1(wireOut[1]), .ctrl(ctrl[0]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_1(.inData_0(wireIn[2]), .inData_1(wireIn[3]), .outData_0(wireOut[2]), .outData_1(wireOut[3]), .ctrl(ctrl[1]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_2(.inData_0(wireIn[4]), .inData_1(wireIn[5]), .outData_0(wireOut[4]), .outData_1(wireOut[5]), .ctrl(ctrl[2]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_3(.inData_0(wireIn[6]), .inData_1(wireIn[7]), .outData_0(wireOut[6]), .outData_1(wireOut[7]), .ctrl(ctrl[3]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_4(.inData_0(wireIn[8]), .inData_1(wireIn[9]), .outData_0(wireOut[8]), .outData_1(wireOut[9]), .ctrl(ctrl[4]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_5(.inData_0(wireIn[10]), .inData_1(wireIn[11]), .outData_0(wireOut[10]), .outData_1(wireOut[11]), .ctrl(ctrl[5]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_6(.inData_0(wireIn[12]), .inData_1(wireIn[13]), .outData_0(wireOut[12]), .outData_1(wireOut[13]), .ctrl(ctrl[6]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_7(.inData_0(wireIn[14]), .inData_1(wireIn[15]), .outData_0(wireOut[14]), .outData_1(wireOut[15]), .ctrl(ctrl[7]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_8(.inData_0(wireIn[16]), .inData_1(wireIn[17]), .outData_0(wireOut[16]), .outData_1(wireOut[17]), .ctrl(ctrl[8]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_9(.inData_0(wireIn[18]), .inData_1(wireIn[19]), .outData_0(wireOut[18]), .outData_1(wireOut[19]), .ctrl(ctrl[9]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_10(.inData_0(wireIn[20]), .inData_1(wireIn[21]), .outData_0(wireOut[20]), .outData_1(wireOut[21]), .ctrl(ctrl[10]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_11(.inData_0(wireIn[22]), .inData_1(wireIn[23]), .outData_0(wireOut[22]), .outData_1(wireOut[23]), .ctrl(ctrl[11]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_12(.inData_0(wireIn[24]), .inData_1(wireIn[25]), .outData_0(wireOut[24]), .outData_1(wireOut[25]), .ctrl(ctrl[12]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_13(.inData_0(wireIn[26]), .inData_1(wireIn[27]), .outData_0(wireOut[26]), .outData_1(wireOut[27]), .ctrl(ctrl[13]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_14(.inData_0(wireIn[28]), .inData_1(wireIn[29]), .outData_0(wireOut[28]), .outData_1(wireOut[29]), .ctrl(ctrl[14]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_15(.inData_0(wireIn[30]), .inData_1(wireIn[31]), .outData_0(wireOut[30]), .outData_1(wireOut[31]), .ctrl(ctrl[15]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_16(.inData_0(wireIn[32]), .inData_1(wireIn[33]), .outData_0(wireOut[32]), .outData_1(wireOut[33]), .ctrl(ctrl[16]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_17(.inData_0(wireIn[34]), .inData_1(wireIn[35]), .outData_0(wireOut[34]), .outData_1(wireOut[35]), .ctrl(ctrl[17]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_18(.inData_0(wireIn[36]), .inData_1(wireIn[37]), .outData_0(wireOut[36]), .outData_1(wireOut[37]), .ctrl(ctrl[18]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_19(.inData_0(wireIn[38]), .inData_1(wireIn[39]), .outData_0(wireOut[38]), .outData_1(wireOut[39]), .ctrl(ctrl[19]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_20(.inData_0(wireIn[40]), .inData_1(wireIn[41]), .outData_0(wireOut[40]), .outData_1(wireOut[41]), .ctrl(ctrl[20]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_21(.inData_0(wireIn[42]), .inData_1(wireIn[43]), .outData_0(wireOut[42]), .outData_1(wireOut[43]), .ctrl(ctrl[21]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_22(.inData_0(wireIn[44]), .inData_1(wireIn[45]), .outData_0(wireOut[44]), .outData_1(wireOut[45]), .ctrl(ctrl[22]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_23(.inData_0(wireIn[46]), .inData_1(wireIn[47]), .outData_0(wireOut[46]), .outData_1(wireOut[47]), .ctrl(ctrl[23]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_24(.inData_0(wireIn[48]), .inData_1(wireIn[49]), .outData_0(wireOut[48]), .outData_1(wireOut[49]), .ctrl(ctrl[24]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_25(.inData_0(wireIn[50]), .inData_1(wireIn[51]), .outData_0(wireOut[50]), .outData_1(wireOut[51]), .ctrl(ctrl[25]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_26(.inData_0(wireIn[52]), .inData_1(wireIn[53]), .outData_0(wireOut[52]), .outData_1(wireOut[53]), .ctrl(ctrl[26]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_27(.inData_0(wireIn[54]), .inData_1(wireIn[55]), .outData_0(wireOut[54]), .outData_1(wireOut[55]), .ctrl(ctrl[27]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_28(.inData_0(wireIn[56]), .inData_1(wireIn[57]), .outData_0(wireOut[56]), .outData_1(wireOut[57]), .ctrl(ctrl[28]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_29(.inData_0(wireIn[58]), .inData_1(wireIn[59]), .outData_0(wireOut[58]), .outData_1(wireOut[59]), .ctrl(ctrl[29]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_30(.inData_0(wireIn[60]), .inData_1(wireIn[61]), .outData_0(wireOut[60]), .outData_1(wireOut[61]), .ctrl(ctrl[30]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_31(.inData_0(wireIn[62]), .inData_1(wireIn[63]), .outData_0(wireOut[62]), .outData_1(wireOut[63]), .ctrl(ctrl[31]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_32(.inData_0(wireIn[64]), .inData_1(wireIn[65]), .outData_0(wireOut[64]), .outData_1(wireOut[65]), .ctrl(ctrl[32]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_33(.inData_0(wireIn[66]), .inData_1(wireIn[67]), .outData_0(wireOut[66]), .outData_1(wireOut[67]), .ctrl(ctrl[33]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_34(.inData_0(wireIn[68]), .inData_1(wireIn[69]), .outData_0(wireOut[68]), .outData_1(wireOut[69]), .ctrl(ctrl[34]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_35(.inData_0(wireIn[70]), .inData_1(wireIn[71]), .outData_0(wireOut[70]), .outData_1(wireOut[71]), .ctrl(ctrl[35]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_36(.inData_0(wireIn[72]), .inData_1(wireIn[73]), .outData_0(wireOut[72]), .outData_1(wireOut[73]), .ctrl(ctrl[36]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_37(.inData_0(wireIn[74]), .inData_1(wireIn[75]), .outData_0(wireOut[74]), .outData_1(wireOut[75]), .ctrl(ctrl[37]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_38(.inData_0(wireIn[76]), .inData_1(wireIn[77]), .outData_0(wireOut[76]), .outData_1(wireOut[77]), .ctrl(ctrl[38]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_39(.inData_0(wireIn[78]), .inData_1(wireIn[79]), .outData_0(wireOut[78]), .outData_1(wireOut[79]), .ctrl(ctrl[39]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_40(.inData_0(wireIn[80]), .inData_1(wireIn[81]), .outData_0(wireOut[80]), .outData_1(wireOut[81]), .ctrl(ctrl[40]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_41(.inData_0(wireIn[82]), .inData_1(wireIn[83]), .outData_0(wireOut[82]), .outData_1(wireOut[83]), .ctrl(ctrl[41]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_42(.inData_0(wireIn[84]), .inData_1(wireIn[85]), .outData_0(wireOut[84]), .outData_1(wireOut[85]), .ctrl(ctrl[42]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_43(.inData_0(wireIn[86]), .inData_1(wireIn[87]), .outData_0(wireOut[86]), .outData_1(wireOut[87]), .ctrl(ctrl[43]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_44(.inData_0(wireIn[88]), .inData_1(wireIn[89]), .outData_0(wireOut[88]), .outData_1(wireOut[89]), .ctrl(ctrl[44]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_45(.inData_0(wireIn[90]), .inData_1(wireIn[91]), .outData_0(wireOut[90]), .outData_1(wireOut[91]), .ctrl(ctrl[45]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_46(.inData_0(wireIn[92]), .inData_1(wireIn[93]), .outData_0(wireOut[92]), .outData_1(wireOut[93]), .ctrl(ctrl[46]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_47(.inData_0(wireIn[94]), .inData_1(wireIn[95]), .outData_0(wireOut[94]), .outData_1(wireOut[95]), .ctrl(ctrl[47]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_48(.inData_0(wireIn[96]), .inData_1(wireIn[97]), .outData_0(wireOut[96]), .outData_1(wireOut[97]), .ctrl(ctrl[48]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_49(.inData_0(wireIn[98]), .inData_1(wireIn[99]), .outData_0(wireOut[98]), .outData_1(wireOut[99]), .ctrl(ctrl[49]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_50(.inData_0(wireIn[100]), .inData_1(wireIn[101]), .outData_0(wireOut[100]), .outData_1(wireOut[101]), .ctrl(ctrl[50]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_51(.inData_0(wireIn[102]), .inData_1(wireIn[103]), .outData_0(wireOut[102]), .outData_1(wireOut[103]), .ctrl(ctrl[51]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_52(.inData_0(wireIn[104]), .inData_1(wireIn[105]), .outData_0(wireOut[104]), .outData_1(wireOut[105]), .ctrl(ctrl[52]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_53(.inData_0(wireIn[106]), .inData_1(wireIn[107]), .outData_0(wireOut[106]), .outData_1(wireOut[107]), .ctrl(ctrl[53]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_54(.inData_0(wireIn[108]), .inData_1(wireIn[109]), .outData_0(wireOut[108]), .outData_1(wireOut[109]), .ctrl(ctrl[54]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_55(.inData_0(wireIn[110]), .inData_1(wireIn[111]), .outData_0(wireOut[110]), .outData_1(wireOut[111]), .ctrl(ctrl[55]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_56(.inData_0(wireIn[112]), .inData_1(wireIn[113]), .outData_0(wireOut[112]), .outData_1(wireOut[113]), .ctrl(ctrl[56]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_57(.inData_0(wireIn[114]), .inData_1(wireIn[115]), .outData_0(wireOut[114]), .outData_1(wireOut[115]), .ctrl(ctrl[57]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_58(.inData_0(wireIn[116]), .inData_1(wireIn[117]), .outData_0(wireOut[116]), .outData_1(wireOut[117]), .ctrl(ctrl[58]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_59(.inData_0(wireIn[118]), .inData_1(wireIn[119]), .outData_0(wireOut[118]), .outData_1(wireOut[119]), .ctrl(ctrl[59]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_60(.inData_0(wireIn[120]), .inData_1(wireIn[121]), .outData_0(wireOut[120]), .outData_1(wireOut[121]), .ctrl(ctrl[60]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_61(.inData_0(wireIn[122]), .inData_1(wireIn[123]), .outData_0(wireOut[122]), .outData_1(wireOut[123]), .ctrl(ctrl[61]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_62(.inData_0(wireIn[124]), .inData_1(wireIn[125]), .outData_0(wireOut[124]), .outData_1(wireOut[125]), .ctrl(ctrl[62]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_63(.inData_0(wireIn[126]), .inData_1(wireIn[127]), .outData_0(wireOut[126]), .outData_1(wireOut[127]), .ctrl(ctrl[63]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_64(.inData_0(wireIn[128]), .inData_1(wireIn[129]), .outData_0(wireOut[128]), .outData_1(wireOut[129]), .ctrl(ctrl[64]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_65(.inData_0(wireIn[130]), .inData_1(wireIn[131]), .outData_0(wireOut[130]), .outData_1(wireOut[131]), .ctrl(ctrl[65]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_66(.inData_0(wireIn[132]), .inData_1(wireIn[133]), .outData_0(wireOut[132]), .outData_1(wireOut[133]), .ctrl(ctrl[66]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_67(.inData_0(wireIn[134]), .inData_1(wireIn[135]), .outData_0(wireOut[134]), .outData_1(wireOut[135]), .ctrl(ctrl[67]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_68(.inData_0(wireIn[136]), .inData_1(wireIn[137]), .outData_0(wireOut[136]), .outData_1(wireOut[137]), .ctrl(ctrl[68]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_69(.inData_0(wireIn[138]), .inData_1(wireIn[139]), .outData_0(wireOut[138]), .outData_1(wireOut[139]), .ctrl(ctrl[69]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_70(.inData_0(wireIn[140]), .inData_1(wireIn[141]), .outData_0(wireOut[140]), .outData_1(wireOut[141]), .ctrl(ctrl[70]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_71(.inData_0(wireIn[142]), .inData_1(wireIn[143]), .outData_0(wireOut[142]), .outData_1(wireOut[143]), .ctrl(ctrl[71]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_72(.inData_0(wireIn[144]), .inData_1(wireIn[145]), .outData_0(wireOut[144]), .outData_1(wireOut[145]), .ctrl(ctrl[72]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_73(.inData_0(wireIn[146]), .inData_1(wireIn[147]), .outData_0(wireOut[146]), .outData_1(wireOut[147]), .ctrl(ctrl[73]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_74(.inData_0(wireIn[148]), .inData_1(wireIn[149]), .outData_0(wireOut[148]), .outData_1(wireOut[149]), .ctrl(ctrl[74]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_75(.inData_0(wireIn[150]), .inData_1(wireIn[151]), .outData_0(wireOut[150]), .outData_1(wireOut[151]), .ctrl(ctrl[75]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_76(.inData_0(wireIn[152]), .inData_1(wireIn[153]), .outData_0(wireOut[152]), .outData_1(wireOut[153]), .ctrl(ctrl[76]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_77(.inData_0(wireIn[154]), .inData_1(wireIn[155]), .outData_0(wireOut[154]), .outData_1(wireOut[155]), .ctrl(ctrl[77]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_78(.inData_0(wireIn[156]), .inData_1(wireIn[157]), .outData_0(wireOut[156]), .outData_1(wireOut[157]), .ctrl(ctrl[78]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_79(.inData_0(wireIn[158]), .inData_1(wireIn[159]), .outData_0(wireOut[158]), .outData_1(wireOut[159]), .ctrl(ctrl[79]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_80(.inData_0(wireIn[160]), .inData_1(wireIn[161]), .outData_0(wireOut[160]), .outData_1(wireOut[161]), .ctrl(ctrl[80]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_81(.inData_0(wireIn[162]), .inData_1(wireIn[163]), .outData_0(wireOut[162]), .outData_1(wireOut[163]), .ctrl(ctrl[81]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_82(.inData_0(wireIn[164]), .inData_1(wireIn[165]), .outData_0(wireOut[164]), .outData_1(wireOut[165]), .ctrl(ctrl[82]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_83(.inData_0(wireIn[166]), .inData_1(wireIn[167]), .outData_0(wireOut[166]), .outData_1(wireOut[167]), .ctrl(ctrl[83]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_84(.inData_0(wireIn[168]), .inData_1(wireIn[169]), .outData_0(wireOut[168]), .outData_1(wireOut[169]), .ctrl(ctrl[84]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_85(.inData_0(wireIn[170]), .inData_1(wireIn[171]), .outData_0(wireOut[170]), .outData_1(wireOut[171]), .ctrl(ctrl[85]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_86(.inData_0(wireIn[172]), .inData_1(wireIn[173]), .outData_0(wireOut[172]), .outData_1(wireOut[173]), .ctrl(ctrl[86]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_87(.inData_0(wireIn[174]), .inData_1(wireIn[175]), .outData_0(wireOut[174]), .outData_1(wireOut[175]), .ctrl(ctrl[87]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_88(.inData_0(wireIn[176]), .inData_1(wireIn[177]), .outData_0(wireOut[176]), .outData_1(wireOut[177]), .ctrl(ctrl[88]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_89(.inData_0(wireIn[178]), .inData_1(wireIn[179]), .outData_0(wireOut[178]), .outData_1(wireOut[179]), .ctrl(ctrl[89]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_90(.inData_0(wireIn[180]), .inData_1(wireIn[181]), .outData_0(wireOut[180]), .outData_1(wireOut[181]), .ctrl(ctrl[90]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_91(.inData_0(wireIn[182]), .inData_1(wireIn[183]), .outData_0(wireOut[182]), .outData_1(wireOut[183]), .ctrl(ctrl[91]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_92(.inData_0(wireIn[184]), .inData_1(wireIn[185]), .outData_0(wireOut[184]), .outData_1(wireOut[185]), .ctrl(ctrl[92]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_93(.inData_0(wireIn[186]), .inData_1(wireIn[187]), .outData_0(wireOut[186]), .outData_1(wireOut[187]), .ctrl(ctrl[93]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_94(.inData_0(wireIn[188]), .inData_1(wireIn[189]), .outData_0(wireOut[188]), .outData_1(wireOut[189]), .ctrl(ctrl[94]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_95(.inData_0(wireIn[190]), .inData_1(wireIn[191]), .outData_0(wireOut[190]), .outData_1(wireOut[191]), .ctrl(ctrl[95]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_96(.inData_0(wireIn[192]), .inData_1(wireIn[193]), .outData_0(wireOut[192]), .outData_1(wireOut[193]), .ctrl(ctrl[96]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_97(.inData_0(wireIn[194]), .inData_1(wireIn[195]), .outData_0(wireOut[194]), .outData_1(wireOut[195]), .ctrl(ctrl[97]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_98(.inData_0(wireIn[196]), .inData_1(wireIn[197]), .outData_0(wireOut[196]), .outData_1(wireOut[197]), .ctrl(ctrl[98]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_99(.inData_0(wireIn[198]), .inData_1(wireIn[199]), .outData_0(wireOut[198]), .outData_1(wireOut[199]), .ctrl(ctrl[99]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_100(.inData_0(wireIn[200]), .inData_1(wireIn[201]), .outData_0(wireOut[200]), .outData_1(wireOut[201]), .ctrl(ctrl[100]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_101(.inData_0(wireIn[202]), .inData_1(wireIn[203]), .outData_0(wireOut[202]), .outData_1(wireOut[203]), .ctrl(ctrl[101]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_102(.inData_0(wireIn[204]), .inData_1(wireIn[205]), .outData_0(wireOut[204]), .outData_1(wireOut[205]), .ctrl(ctrl[102]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_103(.inData_0(wireIn[206]), .inData_1(wireIn[207]), .outData_0(wireOut[206]), .outData_1(wireOut[207]), .ctrl(ctrl[103]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_104(.inData_0(wireIn[208]), .inData_1(wireIn[209]), .outData_0(wireOut[208]), .outData_1(wireOut[209]), .ctrl(ctrl[104]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_105(.inData_0(wireIn[210]), .inData_1(wireIn[211]), .outData_0(wireOut[210]), .outData_1(wireOut[211]), .ctrl(ctrl[105]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_106(.inData_0(wireIn[212]), .inData_1(wireIn[213]), .outData_0(wireOut[212]), .outData_1(wireOut[213]), .ctrl(ctrl[106]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_107(.inData_0(wireIn[214]), .inData_1(wireIn[215]), .outData_0(wireOut[214]), .outData_1(wireOut[215]), .ctrl(ctrl[107]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_108(.inData_0(wireIn[216]), .inData_1(wireIn[217]), .outData_0(wireOut[216]), .outData_1(wireOut[217]), .ctrl(ctrl[108]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_109(.inData_0(wireIn[218]), .inData_1(wireIn[219]), .outData_0(wireOut[218]), .outData_1(wireOut[219]), .ctrl(ctrl[109]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_110(.inData_0(wireIn[220]), .inData_1(wireIn[221]), .outData_0(wireOut[220]), .outData_1(wireOut[221]), .ctrl(ctrl[110]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_111(.inData_0(wireIn[222]), .inData_1(wireIn[223]), .outData_0(wireOut[222]), .outData_1(wireOut[223]), .ctrl(ctrl[111]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_112(.inData_0(wireIn[224]), .inData_1(wireIn[225]), .outData_0(wireOut[224]), .outData_1(wireOut[225]), .ctrl(ctrl[112]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_113(.inData_0(wireIn[226]), .inData_1(wireIn[227]), .outData_0(wireOut[226]), .outData_1(wireOut[227]), .ctrl(ctrl[113]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_114(.inData_0(wireIn[228]), .inData_1(wireIn[229]), .outData_0(wireOut[228]), .outData_1(wireOut[229]), .ctrl(ctrl[114]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_115(.inData_0(wireIn[230]), .inData_1(wireIn[231]), .outData_0(wireOut[230]), .outData_1(wireOut[231]), .ctrl(ctrl[115]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_116(.inData_0(wireIn[232]), .inData_1(wireIn[233]), .outData_0(wireOut[232]), .outData_1(wireOut[233]), .ctrl(ctrl[116]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_117(.inData_0(wireIn[234]), .inData_1(wireIn[235]), .outData_0(wireOut[234]), .outData_1(wireOut[235]), .ctrl(ctrl[117]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_118(.inData_0(wireIn[236]), .inData_1(wireIn[237]), .outData_0(wireOut[236]), .outData_1(wireOut[237]), .ctrl(ctrl[118]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_119(.inData_0(wireIn[238]), .inData_1(wireIn[239]), .outData_0(wireOut[238]), .outData_1(wireOut[239]), .ctrl(ctrl[119]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_120(.inData_0(wireIn[240]), .inData_1(wireIn[241]), .outData_0(wireOut[240]), .outData_1(wireOut[241]), .ctrl(ctrl[120]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_121(.inData_0(wireIn[242]), .inData_1(wireIn[243]), .outData_0(wireOut[242]), .outData_1(wireOut[243]), .ctrl(ctrl[121]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_122(.inData_0(wireIn[244]), .inData_1(wireIn[245]), .outData_0(wireOut[244]), .outData_1(wireOut[245]), .ctrl(ctrl[122]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_123(.inData_0(wireIn[246]), .inData_1(wireIn[247]), .outData_0(wireOut[246]), .outData_1(wireOut[247]), .ctrl(ctrl[123]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_124(.inData_0(wireIn[248]), .inData_1(wireIn[249]), .outData_0(wireOut[248]), .outData_1(wireOut[249]), .ctrl(ctrl[124]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_125(.inData_0(wireIn[250]), .inData_1(wireIn[251]), .outData_0(wireOut[250]), .outData_1(wireOut[251]), .ctrl(ctrl[125]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_126(.inData_0(wireIn[252]), .inData_1(wireIn[253]), .outData_0(wireOut[252]), .outData_1(wireOut[253]), .ctrl(ctrl[126]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_127(.inData_0(wireIn[254]), .inData_1(wireIn[255]), .outData_0(wireOut[254]), .outData_1(wireOut[255]), .ctrl(ctrl[127]), .clk(clk), .rst(rst));
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module wireCon_dp256_st3_R(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  assign wireOut[0] = wireIn[0];    
  assign wireOut[1] = wireIn[16];    
  assign wireOut[2] = wireIn[1];    
  assign wireOut[3] = wireIn[17];    
  assign wireOut[4] = wireIn[2];    
  assign wireOut[5] = wireIn[18];    
  assign wireOut[6] = wireIn[3];    
  assign wireOut[7] = wireIn[19];    
  assign wireOut[8] = wireIn[4];    
  assign wireOut[9] = wireIn[20];    
  assign wireOut[10] = wireIn[5];    
  assign wireOut[11] = wireIn[21];    
  assign wireOut[12] = wireIn[6];    
  assign wireOut[13] = wireIn[22];    
  assign wireOut[14] = wireIn[7];    
  assign wireOut[15] = wireIn[23];    
  assign wireOut[16] = wireIn[8];    
  assign wireOut[17] = wireIn[24];    
  assign wireOut[18] = wireIn[9];    
  assign wireOut[19] = wireIn[25];    
  assign wireOut[20] = wireIn[10];    
  assign wireOut[21] = wireIn[26];    
  assign wireOut[22] = wireIn[11];    
  assign wireOut[23] = wireIn[27];    
  assign wireOut[24] = wireIn[12];    
  assign wireOut[25] = wireIn[28];    
  assign wireOut[26] = wireIn[13];    
  assign wireOut[27] = wireIn[29];    
  assign wireOut[28] = wireIn[14];    
  assign wireOut[29] = wireIn[30];    
  assign wireOut[30] = wireIn[15];    
  assign wireOut[31] = wireIn[31];    
  assign wireOut[32] = wireIn[32];    
  assign wireOut[33] = wireIn[48];    
  assign wireOut[34] = wireIn[33];    
  assign wireOut[35] = wireIn[49];    
  assign wireOut[36] = wireIn[34];    
  assign wireOut[37] = wireIn[50];    
  assign wireOut[38] = wireIn[35];    
  assign wireOut[39] = wireIn[51];    
  assign wireOut[40] = wireIn[36];    
  assign wireOut[41] = wireIn[52];    
  assign wireOut[42] = wireIn[37];    
  assign wireOut[43] = wireIn[53];    
  assign wireOut[44] = wireIn[38];    
  assign wireOut[45] = wireIn[54];    
  assign wireOut[46] = wireIn[39];    
  assign wireOut[47] = wireIn[55];    
  assign wireOut[48] = wireIn[40];    
  assign wireOut[49] = wireIn[56];    
  assign wireOut[50] = wireIn[41];    
  assign wireOut[51] = wireIn[57];    
  assign wireOut[52] = wireIn[42];    
  assign wireOut[53] = wireIn[58];    
  assign wireOut[54] = wireIn[43];    
  assign wireOut[55] = wireIn[59];    
  assign wireOut[56] = wireIn[44];    
  assign wireOut[57] = wireIn[60];    
  assign wireOut[58] = wireIn[45];    
  assign wireOut[59] = wireIn[61];    
  assign wireOut[60] = wireIn[46];    
  assign wireOut[61] = wireIn[62];    
  assign wireOut[62] = wireIn[47];    
  assign wireOut[63] = wireIn[63];    
  assign wireOut[64] = wireIn[64];    
  assign wireOut[65] = wireIn[80];    
  assign wireOut[66] = wireIn[65];    
  assign wireOut[67] = wireIn[81];    
  assign wireOut[68] = wireIn[66];    
  assign wireOut[69] = wireIn[82];    
  assign wireOut[70] = wireIn[67];    
  assign wireOut[71] = wireIn[83];    
  assign wireOut[72] = wireIn[68];    
  assign wireOut[73] = wireIn[84];    
  assign wireOut[74] = wireIn[69];    
  assign wireOut[75] = wireIn[85];    
  assign wireOut[76] = wireIn[70];    
  assign wireOut[77] = wireIn[86];    
  assign wireOut[78] = wireIn[71];    
  assign wireOut[79] = wireIn[87];    
  assign wireOut[80] = wireIn[72];    
  assign wireOut[81] = wireIn[88];    
  assign wireOut[82] = wireIn[73];    
  assign wireOut[83] = wireIn[89];    
  assign wireOut[84] = wireIn[74];    
  assign wireOut[85] = wireIn[90];    
  assign wireOut[86] = wireIn[75];    
  assign wireOut[87] = wireIn[91];    
  assign wireOut[88] = wireIn[76];    
  assign wireOut[89] = wireIn[92];    
  assign wireOut[90] = wireIn[77];    
  assign wireOut[91] = wireIn[93];    
  assign wireOut[92] = wireIn[78];    
  assign wireOut[93] = wireIn[94];    
  assign wireOut[94] = wireIn[79];    
  assign wireOut[95] = wireIn[95];    
  assign wireOut[96] = wireIn[96];    
  assign wireOut[97] = wireIn[112];    
  assign wireOut[98] = wireIn[97];    
  assign wireOut[99] = wireIn[113];    
  assign wireOut[100] = wireIn[98];    
  assign wireOut[101] = wireIn[114];    
  assign wireOut[102] = wireIn[99];    
  assign wireOut[103] = wireIn[115];    
  assign wireOut[104] = wireIn[100];    
  assign wireOut[105] = wireIn[116];    
  assign wireOut[106] = wireIn[101];    
  assign wireOut[107] = wireIn[117];    
  assign wireOut[108] = wireIn[102];    
  assign wireOut[109] = wireIn[118];    
  assign wireOut[110] = wireIn[103];    
  assign wireOut[111] = wireIn[119];    
  assign wireOut[112] = wireIn[104];    
  assign wireOut[113] = wireIn[120];    
  assign wireOut[114] = wireIn[105];    
  assign wireOut[115] = wireIn[121];    
  assign wireOut[116] = wireIn[106];    
  assign wireOut[117] = wireIn[122];    
  assign wireOut[118] = wireIn[107];    
  assign wireOut[119] = wireIn[123];    
  assign wireOut[120] = wireIn[108];    
  assign wireOut[121] = wireIn[124];    
  assign wireOut[122] = wireIn[109];    
  assign wireOut[123] = wireIn[125];    
  assign wireOut[124] = wireIn[110];    
  assign wireOut[125] = wireIn[126];    
  assign wireOut[126] = wireIn[111];    
  assign wireOut[127] = wireIn[127];    
  assign wireOut[128] = wireIn[128];    
  assign wireOut[129] = wireIn[144];    
  assign wireOut[130] = wireIn[129];    
  assign wireOut[131] = wireIn[145];    
  assign wireOut[132] = wireIn[130];    
  assign wireOut[133] = wireIn[146];    
  assign wireOut[134] = wireIn[131];    
  assign wireOut[135] = wireIn[147];    
  assign wireOut[136] = wireIn[132];    
  assign wireOut[137] = wireIn[148];    
  assign wireOut[138] = wireIn[133];    
  assign wireOut[139] = wireIn[149];    
  assign wireOut[140] = wireIn[134];    
  assign wireOut[141] = wireIn[150];    
  assign wireOut[142] = wireIn[135];    
  assign wireOut[143] = wireIn[151];    
  assign wireOut[144] = wireIn[136];    
  assign wireOut[145] = wireIn[152];    
  assign wireOut[146] = wireIn[137];    
  assign wireOut[147] = wireIn[153];    
  assign wireOut[148] = wireIn[138];    
  assign wireOut[149] = wireIn[154];    
  assign wireOut[150] = wireIn[139];    
  assign wireOut[151] = wireIn[155];    
  assign wireOut[152] = wireIn[140];    
  assign wireOut[153] = wireIn[156];    
  assign wireOut[154] = wireIn[141];    
  assign wireOut[155] = wireIn[157];    
  assign wireOut[156] = wireIn[142];    
  assign wireOut[157] = wireIn[158];    
  assign wireOut[158] = wireIn[143];    
  assign wireOut[159] = wireIn[159];    
  assign wireOut[160] = wireIn[160];    
  assign wireOut[161] = wireIn[176];    
  assign wireOut[162] = wireIn[161];    
  assign wireOut[163] = wireIn[177];    
  assign wireOut[164] = wireIn[162];    
  assign wireOut[165] = wireIn[178];    
  assign wireOut[166] = wireIn[163];    
  assign wireOut[167] = wireIn[179];    
  assign wireOut[168] = wireIn[164];    
  assign wireOut[169] = wireIn[180];    
  assign wireOut[170] = wireIn[165];    
  assign wireOut[171] = wireIn[181];    
  assign wireOut[172] = wireIn[166];    
  assign wireOut[173] = wireIn[182];    
  assign wireOut[174] = wireIn[167];    
  assign wireOut[175] = wireIn[183];    
  assign wireOut[176] = wireIn[168];    
  assign wireOut[177] = wireIn[184];    
  assign wireOut[178] = wireIn[169];    
  assign wireOut[179] = wireIn[185];    
  assign wireOut[180] = wireIn[170];    
  assign wireOut[181] = wireIn[186];    
  assign wireOut[182] = wireIn[171];    
  assign wireOut[183] = wireIn[187];    
  assign wireOut[184] = wireIn[172];    
  assign wireOut[185] = wireIn[188];    
  assign wireOut[186] = wireIn[173];    
  assign wireOut[187] = wireIn[189];    
  assign wireOut[188] = wireIn[174];    
  assign wireOut[189] = wireIn[190];    
  assign wireOut[190] = wireIn[175];    
  assign wireOut[191] = wireIn[191];    
  assign wireOut[192] = wireIn[192];    
  assign wireOut[193] = wireIn[208];    
  assign wireOut[194] = wireIn[193];    
  assign wireOut[195] = wireIn[209];    
  assign wireOut[196] = wireIn[194];    
  assign wireOut[197] = wireIn[210];    
  assign wireOut[198] = wireIn[195];    
  assign wireOut[199] = wireIn[211];    
  assign wireOut[200] = wireIn[196];    
  assign wireOut[201] = wireIn[212];    
  assign wireOut[202] = wireIn[197];    
  assign wireOut[203] = wireIn[213];    
  assign wireOut[204] = wireIn[198];    
  assign wireOut[205] = wireIn[214];    
  assign wireOut[206] = wireIn[199];    
  assign wireOut[207] = wireIn[215];    
  assign wireOut[208] = wireIn[200];    
  assign wireOut[209] = wireIn[216];    
  assign wireOut[210] = wireIn[201];    
  assign wireOut[211] = wireIn[217];    
  assign wireOut[212] = wireIn[202];    
  assign wireOut[213] = wireIn[218];    
  assign wireOut[214] = wireIn[203];    
  assign wireOut[215] = wireIn[219];    
  assign wireOut[216] = wireIn[204];    
  assign wireOut[217] = wireIn[220];    
  assign wireOut[218] = wireIn[205];    
  assign wireOut[219] = wireIn[221];    
  assign wireOut[220] = wireIn[206];    
  assign wireOut[221] = wireIn[222];    
  assign wireOut[222] = wireIn[207];    
  assign wireOut[223] = wireIn[223];    
  assign wireOut[224] = wireIn[224];    
  assign wireOut[225] = wireIn[240];    
  assign wireOut[226] = wireIn[225];    
  assign wireOut[227] = wireIn[241];    
  assign wireOut[228] = wireIn[226];    
  assign wireOut[229] = wireIn[242];    
  assign wireOut[230] = wireIn[227];    
  assign wireOut[231] = wireIn[243];    
  assign wireOut[232] = wireIn[228];    
  assign wireOut[233] = wireIn[244];    
  assign wireOut[234] = wireIn[229];    
  assign wireOut[235] = wireIn[245];    
  assign wireOut[236] = wireIn[230];    
  assign wireOut[237] = wireIn[246];    
  assign wireOut[238] = wireIn[231];    
  assign wireOut[239] = wireIn[247];    
  assign wireOut[240] = wireIn[232];    
  assign wireOut[241] = wireIn[248];    
  assign wireOut[242] = wireIn[233];    
  assign wireOut[243] = wireIn[249];    
  assign wireOut[244] = wireIn[234];    
  assign wireOut[245] = wireIn[250];    
  assign wireOut[246] = wireIn[235];    
  assign wireOut[247] = wireIn[251];    
  assign wireOut[248] = wireIn[236];    
  assign wireOut[249] = wireIn[252];    
  assign wireOut[250] = wireIn[237];    
  assign wireOut[251] = wireIn[253];    
  assign wireOut[252] = wireIn[238];    
  assign wireOut[253] = wireIn[254];    
  assign wireOut[254] = wireIn[239];    
  assign wireOut[255] = wireIn[255];    
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module switches_stage_st4_0_R(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
ctrl,                            
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;                   
  input [128-1:0] ctrl;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  switch_2_2 switch_inst_0(.inData_0(wireIn[0]), .inData_1(wireIn[1]), .outData_0(wireOut[0]), .outData_1(wireOut[1]), .ctrl(ctrl[0]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_1(.inData_0(wireIn[2]), .inData_1(wireIn[3]), .outData_0(wireOut[2]), .outData_1(wireOut[3]), .ctrl(ctrl[1]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_2(.inData_0(wireIn[4]), .inData_1(wireIn[5]), .outData_0(wireOut[4]), .outData_1(wireOut[5]), .ctrl(ctrl[2]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_3(.inData_0(wireIn[6]), .inData_1(wireIn[7]), .outData_0(wireOut[6]), .outData_1(wireOut[7]), .ctrl(ctrl[3]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_4(.inData_0(wireIn[8]), .inData_1(wireIn[9]), .outData_0(wireOut[8]), .outData_1(wireOut[9]), .ctrl(ctrl[4]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_5(.inData_0(wireIn[10]), .inData_1(wireIn[11]), .outData_0(wireOut[10]), .outData_1(wireOut[11]), .ctrl(ctrl[5]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_6(.inData_0(wireIn[12]), .inData_1(wireIn[13]), .outData_0(wireOut[12]), .outData_1(wireOut[13]), .ctrl(ctrl[6]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_7(.inData_0(wireIn[14]), .inData_1(wireIn[15]), .outData_0(wireOut[14]), .outData_1(wireOut[15]), .ctrl(ctrl[7]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_8(.inData_0(wireIn[16]), .inData_1(wireIn[17]), .outData_0(wireOut[16]), .outData_1(wireOut[17]), .ctrl(ctrl[8]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_9(.inData_0(wireIn[18]), .inData_1(wireIn[19]), .outData_0(wireOut[18]), .outData_1(wireOut[19]), .ctrl(ctrl[9]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_10(.inData_0(wireIn[20]), .inData_1(wireIn[21]), .outData_0(wireOut[20]), .outData_1(wireOut[21]), .ctrl(ctrl[10]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_11(.inData_0(wireIn[22]), .inData_1(wireIn[23]), .outData_0(wireOut[22]), .outData_1(wireOut[23]), .ctrl(ctrl[11]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_12(.inData_0(wireIn[24]), .inData_1(wireIn[25]), .outData_0(wireOut[24]), .outData_1(wireOut[25]), .ctrl(ctrl[12]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_13(.inData_0(wireIn[26]), .inData_1(wireIn[27]), .outData_0(wireOut[26]), .outData_1(wireOut[27]), .ctrl(ctrl[13]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_14(.inData_0(wireIn[28]), .inData_1(wireIn[29]), .outData_0(wireOut[28]), .outData_1(wireOut[29]), .ctrl(ctrl[14]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_15(.inData_0(wireIn[30]), .inData_1(wireIn[31]), .outData_0(wireOut[30]), .outData_1(wireOut[31]), .ctrl(ctrl[15]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_16(.inData_0(wireIn[32]), .inData_1(wireIn[33]), .outData_0(wireOut[32]), .outData_1(wireOut[33]), .ctrl(ctrl[16]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_17(.inData_0(wireIn[34]), .inData_1(wireIn[35]), .outData_0(wireOut[34]), .outData_1(wireOut[35]), .ctrl(ctrl[17]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_18(.inData_0(wireIn[36]), .inData_1(wireIn[37]), .outData_0(wireOut[36]), .outData_1(wireOut[37]), .ctrl(ctrl[18]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_19(.inData_0(wireIn[38]), .inData_1(wireIn[39]), .outData_0(wireOut[38]), .outData_1(wireOut[39]), .ctrl(ctrl[19]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_20(.inData_0(wireIn[40]), .inData_1(wireIn[41]), .outData_0(wireOut[40]), .outData_1(wireOut[41]), .ctrl(ctrl[20]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_21(.inData_0(wireIn[42]), .inData_1(wireIn[43]), .outData_0(wireOut[42]), .outData_1(wireOut[43]), .ctrl(ctrl[21]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_22(.inData_0(wireIn[44]), .inData_1(wireIn[45]), .outData_0(wireOut[44]), .outData_1(wireOut[45]), .ctrl(ctrl[22]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_23(.inData_0(wireIn[46]), .inData_1(wireIn[47]), .outData_0(wireOut[46]), .outData_1(wireOut[47]), .ctrl(ctrl[23]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_24(.inData_0(wireIn[48]), .inData_1(wireIn[49]), .outData_0(wireOut[48]), .outData_1(wireOut[49]), .ctrl(ctrl[24]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_25(.inData_0(wireIn[50]), .inData_1(wireIn[51]), .outData_0(wireOut[50]), .outData_1(wireOut[51]), .ctrl(ctrl[25]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_26(.inData_0(wireIn[52]), .inData_1(wireIn[53]), .outData_0(wireOut[52]), .outData_1(wireOut[53]), .ctrl(ctrl[26]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_27(.inData_0(wireIn[54]), .inData_1(wireIn[55]), .outData_0(wireOut[54]), .outData_1(wireOut[55]), .ctrl(ctrl[27]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_28(.inData_0(wireIn[56]), .inData_1(wireIn[57]), .outData_0(wireOut[56]), .outData_1(wireOut[57]), .ctrl(ctrl[28]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_29(.inData_0(wireIn[58]), .inData_1(wireIn[59]), .outData_0(wireOut[58]), .outData_1(wireOut[59]), .ctrl(ctrl[29]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_30(.inData_0(wireIn[60]), .inData_1(wireIn[61]), .outData_0(wireOut[60]), .outData_1(wireOut[61]), .ctrl(ctrl[30]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_31(.inData_0(wireIn[62]), .inData_1(wireIn[63]), .outData_0(wireOut[62]), .outData_1(wireOut[63]), .ctrl(ctrl[31]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_32(.inData_0(wireIn[64]), .inData_1(wireIn[65]), .outData_0(wireOut[64]), .outData_1(wireOut[65]), .ctrl(ctrl[32]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_33(.inData_0(wireIn[66]), .inData_1(wireIn[67]), .outData_0(wireOut[66]), .outData_1(wireOut[67]), .ctrl(ctrl[33]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_34(.inData_0(wireIn[68]), .inData_1(wireIn[69]), .outData_0(wireOut[68]), .outData_1(wireOut[69]), .ctrl(ctrl[34]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_35(.inData_0(wireIn[70]), .inData_1(wireIn[71]), .outData_0(wireOut[70]), .outData_1(wireOut[71]), .ctrl(ctrl[35]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_36(.inData_0(wireIn[72]), .inData_1(wireIn[73]), .outData_0(wireOut[72]), .outData_1(wireOut[73]), .ctrl(ctrl[36]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_37(.inData_0(wireIn[74]), .inData_1(wireIn[75]), .outData_0(wireOut[74]), .outData_1(wireOut[75]), .ctrl(ctrl[37]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_38(.inData_0(wireIn[76]), .inData_1(wireIn[77]), .outData_0(wireOut[76]), .outData_1(wireOut[77]), .ctrl(ctrl[38]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_39(.inData_0(wireIn[78]), .inData_1(wireIn[79]), .outData_0(wireOut[78]), .outData_1(wireOut[79]), .ctrl(ctrl[39]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_40(.inData_0(wireIn[80]), .inData_1(wireIn[81]), .outData_0(wireOut[80]), .outData_1(wireOut[81]), .ctrl(ctrl[40]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_41(.inData_0(wireIn[82]), .inData_1(wireIn[83]), .outData_0(wireOut[82]), .outData_1(wireOut[83]), .ctrl(ctrl[41]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_42(.inData_0(wireIn[84]), .inData_1(wireIn[85]), .outData_0(wireOut[84]), .outData_1(wireOut[85]), .ctrl(ctrl[42]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_43(.inData_0(wireIn[86]), .inData_1(wireIn[87]), .outData_0(wireOut[86]), .outData_1(wireOut[87]), .ctrl(ctrl[43]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_44(.inData_0(wireIn[88]), .inData_1(wireIn[89]), .outData_0(wireOut[88]), .outData_1(wireOut[89]), .ctrl(ctrl[44]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_45(.inData_0(wireIn[90]), .inData_1(wireIn[91]), .outData_0(wireOut[90]), .outData_1(wireOut[91]), .ctrl(ctrl[45]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_46(.inData_0(wireIn[92]), .inData_1(wireIn[93]), .outData_0(wireOut[92]), .outData_1(wireOut[93]), .ctrl(ctrl[46]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_47(.inData_0(wireIn[94]), .inData_1(wireIn[95]), .outData_0(wireOut[94]), .outData_1(wireOut[95]), .ctrl(ctrl[47]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_48(.inData_0(wireIn[96]), .inData_1(wireIn[97]), .outData_0(wireOut[96]), .outData_1(wireOut[97]), .ctrl(ctrl[48]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_49(.inData_0(wireIn[98]), .inData_1(wireIn[99]), .outData_0(wireOut[98]), .outData_1(wireOut[99]), .ctrl(ctrl[49]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_50(.inData_0(wireIn[100]), .inData_1(wireIn[101]), .outData_0(wireOut[100]), .outData_1(wireOut[101]), .ctrl(ctrl[50]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_51(.inData_0(wireIn[102]), .inData_1(wireIn[103]), .outData_0(wireOut[102]), .outData_1(wireOut[103]), .ctrl(ctrl[51]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_52(.inData_0(wireIn[104]), .inData_1(wireIn[105]), .outData_0(wireOut[104]), .outData_1(wireOut[105]), .ctrl(ctrl[52]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_53(.inData_0(wireIn[106]), .inData_1(wireIn[107]), .outData_0(wireOut[106]), .outData_1(wireOut[107]), .ctrl(ctrl[53]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_54(.inData_0(wireIn[108]), .inData_1(wireIn[109]), .outData_0(wireOut[108]), .outData_1(wireOut[109]), .ctrl(ctrl[54]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_55(.inData_0(wireIn[110]), .inData_1(wireIn[111]), .outData_0(wireOut[110]), .outData_1(wireOut[111]), .ctrl(ctrl[55]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_56(.inData_0(wireIn[112]), .inData_1(wireIn[113]), .outData_0(wireOut[112]), .outData_1(wireOut[113]), .ctrl(ctrl[56]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_57(.inData_0(wireIn[114]), .inData_1(wireIn[115]), .outData_0(wireOut[114]), .outData_1(wireOut[115]), .ctrl(ctrl[57]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_58(.inData_0(wireIn[116]), .inData_1(wireIn[117]), .outData_0(wireOut[116]), .outData_1(wireOut[117]), .ctrl(ctrl[58]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_59(.inData_0(wireIn[118]), .inData_1(wireIn[119]), .outData_0(wireOut[118]), .outData_1(wireOut[119]), .ctrl(ctrl[59]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_60(.inData_0(wireIn[120]), .inData_1(wireIn[121]), .outData_0(wireOut[120]), .outData_1(wireOut[121]), .ctrl(ctrl[60]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_61(.inData_0(wireIn[122]), .inData_1(wireIn[123]), .outData_0(wireOut[122]), .outData_1(wireOut[123]), .ctrl(ctrl[61]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_62(.inData_0(wireIn[124]), .inData_1(wireIn[125]), .outData_0(wireOut[124]), .outData_1(wireOut[125]), .ctrl(ctrl[62]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_63(.inData_0(wireIn[126]), .inData_1(wireIn[127]), .outData_0(wireOut[126]), .outData_1(wireOut[127]), .ctrl(ctrl[63]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_64(.inData_0(wireIn[128]), .inData_1(wireIn[129]), .outData_0(wireOut[128]), .outData_1(wireOut[129]), .ctrl(ctrl[64]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_65(.inData_0(wireIn[130]), .inData_1(wireIn[131]), .outData_0(wireOut[130]), .outData_1(wireOut[131]), .ctrl(ctrl[65]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_66(.inData_0(wireIn[132]), .inData_1(wireIn[133]), .outData_0(wireOut[132]), .outData_1(wireOut[133]), .ctrl(ctrl[66]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_67(.inData_0(wireIn[134]), .inData_1(wireIn[135]), .outData_0(wireOut[134]), .outData_1(wireOut[135]), .ctrl(ctrl[67]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_68(.inData_0(wireIn[136]), .inData_1(wireIn[137]), .outData_0(wireOut[136]), .outData_1(wireOut[137]), .ctrl(ctrl[68]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_69(.inData_0(wireIn[138]), .inData_1(wireIn[139]), .outData_0(wireOut[138]), .outData_1(wireOut[139]), .ctrl(ctrl[69]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_70(.inData_0(wireIn[140]), .inData_1(wireIn[141]), .outData_0(wireOut[140]), .outData_1(wireOut[141]), .ctrl(ctrl[70]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_71(.inData_0(wireIn[142]), .inData_1(wireIn[143]), .outData_0(wireOut[142]), .outData_1(wireOut[143]), .ctrl(ctrl[71]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_72(.inData_0(wireIn[144]), .inData_1(wireIn[145]), .outData_0(wireOut[144]), .outData_1(wireOut[145]), .ctrl(ctrl[72]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_73(.inData_0(wireIn[146]), .inData_1(wireIn[147]), .outData_0(wireOut[146]), .outData_1(wireOut[147]), .ctrl(ctrl[73]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_74(.inData_0(wireIn[148]), .inData_1(wireIn[149]), .outData_0(wireOut[148]), .outData_1(wireOut[149]), .ctrl(ctrl[74]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_75(.inData_0(wireIn[150]), .inData_1(wireIn[151]), .outData_0(wireOut[150]), .outData_1(wireOut[151]), .ctrl(ctrl[75]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_76(.inData_0(wireIn[152]), .inData_1(wireIn[153]), .outData_0(wireOut[152]), .outData_1(wireOut[153]), .ctrl(ctrl[76]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_77(.inData_0(wireIn[154]), .inData_1(wireIn[155]), .outData_0(wireOut[154]), .outData_1(wireOut[155]), .ctrl(ctrl[77]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_78(.inData_0(wireIn[156]), .inData_1(wireIn[157]), .outData_0(wireOut[156]), .outData_1(wireOut[157]), .ctrl(ctrl[78]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_79(.inData_0(wireIn[158]), .inData_1(wireIn[159]), .outData_0(wireOut[158]), .outData_1(wireOut[159]), .ctrl(ctrl[79]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_80(.inData_0(wireIn[160]), .inData_1(wireIn[161]), .outData_0(wireOut[160]), .outData_1(wireOut[161]), .ctrl(ctrl[80]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_81(.inData_0(wireIn[162]), .inData_1(wireIn[163]), .outData_0(wireOut[162]), .outData_1(wireOut[163]), .ctrl(ctrl[81]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_82(.inData_0(wireIn[164]), .inData_1(wireIn[165]), .outData_0(wireOut[164]), .outData_1(wireOut[165]), .ctrl(ctrl[82]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_83(.inData_0(wireIn[166]), .inData_1(wireIn[167]), .outData_0(wireOut[166]), .outData_1(wireOut[167]), .ctrl(ctrl[83]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_84(.inData_0(wireIn[168]), .inData_1(wireIn[169]), .outData_0(wireOut[168]), .outData_1(wireOut[169]), .ctrl(ctrl[84]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_85(.inData_0(wireIn[170]), .inData_1(wireIn[171]), .outData_0(wireOut[170]), .outData_1(wireOut[171]), .ctrl(ctrl[85]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_86(.inData_0(wireIn[172]), .inData_1(wireIn[173]), .outData_0(wireOut[172]), .outData_1(wireOut[173]), .ctrl(ctrl[86]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_87(.inData_0(wireIn[174]), .inData_1(wireIn[175]), .outData_0(wireOut[174]), .outData_1(wireOut[175]), .ctrl(ctrl[87]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_88(.inData_0(wireIn[176]), .inData_1(wireIn[177]), .outData_0(wireOut[176]), .outData_1(wireOut[177]), .ctrl(ctrl[88]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_89(.inData_0(wireIn[178]), .inData_1(wireIn[179]), .outData_0(wireOut[178]), .outData_1(wireOut[179]), .ctrl(ctrl[89]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_90(.inData_0(wireIn[180]), .inData_1(wireIn[181]), .outData_0(wireOut[180]), .outData_1(wireOut[181]), .ctrl(ctrl[90]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_91(.inData_0(wireIn[182]), .inData_1(wireIn[183]), .outData_0(wireOut[182]), .outData_1(wireOut[183]), .ctrl(ctrl[91]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_92(.inData_0(wireIn[184]), .inData_1(wireIn[185]), .outData_0(wireOut[184]), .outData_1(wireOut[185]), .ctrl(ctrl[92]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_93(.inData_0(wireIn[186]), .inData_1(wireIn[187]), .outData_0(wireOut[186]), .outData_1(wireOut[187]), .ctrl(ctrl[93]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_94(.inData_0(wireIn[188]), .inData_1(wireIn[189]), .outData_0(wireOut[188]), .outData_1(wireOut[189]), .ctrl(ctrl[94]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_95(.inData_0(wireIn[190]), .inData_1(wireIn[191]), .outData_0(wireOut[190]), .outData_1(wireOut[191]), .ctrl(ctrl[95]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_96(.inData_0(wireIn[192]), .inData_1(wireIn[193]), .outData_0(wireOut[192]), .outData_1(wireOut[193]), .ctrl(ctrl[96]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_97(.inData_0(wireIn[194]), .inData_1(wireIn[195]), .outData_0(wireOut[194]), .outData_1(wireOut[195]), .ctrl(ctrl[97]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_98(.inData_0(wireIn[196]), .inData_1(wireIn[197]), .outData_0(wireOut[196]), .outData_1(wireOut[197]), .ctrl(ctrl[98]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_99(.inData_0(wireIn[198]), .inData_1(wireIn[199]), .outData_0(wireOut[198]), .outData_1(wireOut[199]), .ctrl(ctrl[99]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_100(.inData_0(wireIn[200]), .inData_1(wireIn[201]), .outData_0(wireOut[200]), .outData_1(wireOut[201]), .ctrl(ctrl[100]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_101(.inData_0(wireIn[202]), .inData_1(wireIn[203]), .outData_0(wireOut[202]), .outData_1(wireOut[203]), .ctrl(ctrl[101]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_102(.inData_0(wireIn[204]), .inData_1(wireIn[205]), .outData_0(wireOut[204]), .outData_1(wireOut[205]), .ctrl(ctrl[102]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_103(.inData_0(wireIn[206]), .inData_1(wireIn[207]), .outData_0(wireOut[206]), .outData_1(wireOut[207]), .ctrl(ctrl[103]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_104(.inData_0(wireIn[208]), .inData_1(wireIn[209]), .outData_0(wireOut[208]), .outData_1(wireOut[209]), .ctrl(ctrl[104]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_105(.inData_0(wireIn[210]), .inData_1(wireIn[211]), .outData_0(wireOut[210]), .outData_1(wireOut[211]), .ctrl(ctrl[105]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_106(.inData_0(wireIn[212]), .inData_1(wireIn[213]), .outData_0(wireOut[212]), .outData_1(wireOut[213]), .ctrl(ctrl[106]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_107(.inData_0(wireIn[214]), .inData_1(wireIn[215]), .outData_0(wireOut[214]), .outData_1(wireOut[215]), .ctrl(ctrl[107]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_108(.inData_0(wireIn[216]), .inData_1(wireIn[217]), .outData_0(wireOut[216]), .outData_1(wireOut[217]), .ctrl(ctrl[108]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_109(.inData_0(wireIn[218]), .inData_1(wireIn[219]), .outData_0(wireOut[218]), .outData_1(wireOut[219]), .ctrl(ctrl[109]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_110(.inData_0(wireIn[220]), .inData_1(wireIn[221]), .outData_0(wireOut[220]), .outData_1(wireOut[221]), .ctrl(ctrl[110]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_111(.inData_0(wireIn[222]), .inData_1(wireIn[223]), .outData_0(wireOut[222]), .outData_1(wireOut[223]), .ctrl(ctrl[111]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_112(.inData_0(wireIn[224]), .inData_1(wireIn[225]), .outData_0(wireOut[224]), .outData_1(wireOut[225]), .ctrl(ctrl[112]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_113(.inData_0(wireIn[226]), .inData_1(wireIn[227]), .outData_0(wireOut[226]), .outData_1(wireOut[227]), .ctrl(ctrl[113]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_114(.inData_0(wireIn[228]), .inData_1(wireIn[229]), .outData_0(wireOut[228]), .outData_1(wireOut[229]), .ctrl(ctrl[114]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_115(.inData_0(wireIn[230]), .inData_1(wireIn[231]), .outData_0(wireOut[230]), .outData_1(wireOut[231]), .ctrl(ctrl[115]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_116(.inData_0(wireIn[232]), .inData_1(wireIn[233]), .outData_0(wireOut[232]), .outData_1(wireOut[233]), .ctrl(ctrl[116]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_117(.inData_0(wireIn[234]), .inData_1(wireIn[235]), .outData_0(wireOut[234]), .outData_1(wireOut[235]), .ctrl(ctrl[117]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_118(.inData_0(wireIn[236]), .inData_1(wireIn[237]), .outData_0(wireOut[236]), .outData_1(wireOut[237]), .ctrl(ctrl[118]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_119(.inData_0(wireIn[238]), .inData_1(wireIn[239]), .outData_0(wireOut[238]), .outData_1(wireOut[239]), .ctrl(ctrl[119]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_120(.inData_0(wireIn[240]), .inData_1(wireIn[241]), .outData_0(wireOut[240]), .outData_1(wireOut[241]), .ctrl(ctrl[120]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_121(.inData_0(wireIn[242]), .inData_1(wireIn[243]), .outData_0(wireOut[242]), .outData_1(wireOut[243]), .ctrl(ctrl[121]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_122(.inData_0(wireIn[244]), .inData_1(wireIn[245]), .outData_0(wireOut[244]), .outData_1(wireOut[245]), .ctrl(ctrl[122]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_123(.inData_0(wireIn[246]), .inData_1(wireIn[247]), .outData_0(wireOut[246]), .outData_1(wireOut[247]), .ctrl(ctrl[123]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_124(.inData_0(wireIn[248]), .inData_1(wireIn[249]), .outData_0(wireOut[248]), .outData_1(wireOut[249]), .ctrl(ctrl[124]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_125(.inData_0(wireIn[250]), .inData_1(wireIn[251]), .outData_0(wireOut[250]), .outData_1(wireOut[251]), .ctrl(ctrl[125]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_126(.inData_0(wireIn[252]), .inData_1(wireIn[253]), .outData_0(wireOut[252]), .outData_1(wireOut[253]), .ctrl(ctrl[126]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_127(.inData_0(wireIn[254]), .inData_1(wireIn[255]), .outData_0(wireOut[254]), .outData_1(wireOut[255]), .ctrl(ctrl[127]), .clk(clk), .rst(rst));
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module wireCon_dp256_st4_R(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  assign wireOut[0] = wireIn[0];    
  assign wireOut[1] = wireIn[8];    
  assign wireOut[2] = wireIn[1];    
  assign wireOut[3] = wireIn[9];    
  assign wireOut[4] = wireIn[2];    
  assign wireOut[5] = wireIn[10];    
  assign wireOut[6] = wireIn[3];    
  assign wireOut[7] = wireIn[11];    
  assign wireOut[8] = wireIn[4];    
  assign wireOut[9] = wireIn[12];    
  assign wireOut[10] = wireIn[5];    
  assign wireOut[11] = wireIn[13];    
  assign wireOut[12] = wireIn[6];    
  assign wireOut[13] = wireIn[14];    
  assign wireOut[14] = wireIn[7];    
  assign wireOut[15] = wireIn[15];    
  assign wireOut[16] = wireIn[16];    
  assign wireOut[17] = wireIn[24];    
  assign wireOut[18] = wireIn[17];    
  assign wireOut[19] = wireIn[25];    
  assign wireOut[20] = wireIn[18];    
  assign wireOut[21] = wireIn[26];    
  assign wireOut[22] = wireIn[19];    
  assign wireOut[23] = wireIn[27];    
  assign wireOut[24] = wireIn[20];    
  assign wireOut[25] = wireIn[28];    
  assign wireOut[26] = wireIn[21];    
  assign wireOut[27] = wireIn[29];    
  assign wireOut[28] = wireIn[22];    
  assign wireOut[29] = wireIn[30];    
  assign wireOut[30] = wireIn[23];    
  assign wireOut[31] = wireIn[31];    
  assign wireOut[32] = wireIn[32];    
  assign wireOut[33] = wireIn[40];    
  assign wireOut[34] = wireIn[33];    
  assign wireOut[35] = wireIn[41];    
  assign wireOut[36] = wireIn[34];    
  assign wireOut[37] = wireIn[42];    
  assign wireOut[38] = wireIn[35];    
  assign wireOut[39] = wireIn[43];    
  assign wireOut[40] = wireIn[36];    
  assign wireOut[41] = wireIn[44];    
  assign wireOut[42] = wireIn[37];    
  assign wireOut[43] = wireIn[45];    
  assign wireOut[44] = wireIn[38];    
  assign wireOut[45] = wireIn[46];    
  assign wireOut[46] = wireIn[39];    
  assign wireOut[47] = wireIn[47];    
  assign wireOut[48] = wireIn[48];    
  assign wireOut[49] = wireIn[56];    
  assign wireOut[50] = wireIn[49];    
  assign wireOut[51] = wireIn[57];    
  assign wireOut[52] = wireIn[50];    
  assign wireOut[53] = wireIn[58];    
  assign wireOut[54] = wireIn[51];    
  assign wireOut[55] = wireIn[59];    
  assign wireOut[56] = wireIn[52];    
  assign wireOut[57] = wireIn[60];    
  assign wireOut[58] = wireIn[53];    
  assign wireOut[59] = wireIn[61];    
  assign wireOut[60] = wireIn[54];    
  assign wireOut[61] = wireIn[62];    
  assign wireOut[62] = wireIn[55];    
  assign wireOut[63] = wireIn[63];    
  assign wireOut[64] = wireIn[64];    
  assign wireOut[65] = wireIn[72];    
  assign wireOut[66] = wireIn[65];    
  assign wireOut[67] = wireIn[73];    
  assign wireOut[68] = wireIn[66];    
  assign wireOut[69] = wireIn[74];    
  assign wireOut[70] = wireIn[67];    
  assign wireOut[71] = wireIn[75];    
  assign wireOut[72] = wireIn[68];    
  assign wireOut[73] = wireIn[76];    
  assign wireOut[74] = wireIn[69];    
  assign wireOut[75] = wireIn[77];    
  assign wireOut[76] = wireIn[70];    
  assign wireOut[77] = wireIn[78];    
  assign wireOut[78] = wireIn[71];    
  assign wireOut[79] = wireIn[79];    
  assign wireOut[80] = wireIn[80];    
  assign wireOut[81] = wireIn[88];    
  assign wireOut[82] = wireIn[81];    
  assign wireOut[83] = wireIn[89];    
  assign wireOut[84] = wireIn[82];    
  assign wireOut[85] = wireIn[90];    
  assign wireOut[86] = wireIn[83];    
  assign wireOut[87] = wireIn[91];    
  assign wireOut[88] = wireIn[84];    
  assign wireOut[89] = wireIn[92];    
  assign wireOut[90] = wireIn[85];    
  assign wireOut[91] = wireIn[93];    
  assign wireOut[92] = wireIn[86];    
  assign wireOut[93] = wireIn[94];    
  assign wireOut[94] = wireIn[87];    
  assign wireOut[95] = wireIn[95];    
  assign wireOut[96] = wireIn[96];    
  assign wireOut[97] = wireIn[104];    
  assign wireOut[98] = wireIn[97];    
  assign wireOut[99] = wireIn[105];    
  assign wireOut[100] = wireIn[98];    
  assign wireOut[101] = wireIn[106];    
  assign wireOut[102] = wireIn[99];    
  assign wireOut[103] = wireIn[107];    
  assign wireOut[104] = wireIn[100];    
  assign wireOut[105] = wireIn[108];    
  assign wireOut[106] = wireIn[101];    
  assign wireOut[107] = wireIn[109];    
  assign wireOut[108] = wireIn[102];    
  assign wireOut[109] = wireIn[110];    
  assign wireOut[110] = wireIn[103];    
  assign wireOut[111] = wireIn[111];    
  assign wireOut[112] = wireIn[112];    
  assign wireOut[113] = wireIn[120];    
  assign wireOut[114] = wireIn[113];    
  assign wireOut[115] = wireIn[121];    
  assign wireOut[116] = wireIn[114];    
  assign wireOut[117] = wireIn[122];    
  assign wireOut[118] = wireIn[115];    
  assign wireOut[119] = wireIn[123];    
  assign wireOut[120] = wireIn[116];    
  assign wireOut[121] = wireIn[124];    
  assign wireOut[122] = wireIn[117];    
  assign wireOut[123] = wireIn[125];    
  assign wireOut[124] = wireIn[118];    
  assign wireOut[125] = wireIn[126];    
  assign wireOut[126] = wireIn[119];    
  assign wireOut[127] = wireIn[127];    
  assign wireOut[128] = wireIn[128];    
  assign wireOut[129] = wireIn[136];    
  assign wireOut[130] = wireIn[129];    
  assign wireOut[131] = wireIn[137];    
  assign wireOut[132] = wireIn[130];    
  assign wireOut[133] = wireIn[138];    
  assign wireOut[134] = wireIn[131];    
  assign wireOut[135] = wireIn[139];    
  assign wireOut[136] = wireIn[132];    
  assign wireOut[137] = wireIn[140];    
  assign wireOut[138] = wireIn[133];    
  assign wireOut[139] = wireIn[141];    
  assign wireOut[140] = wireIn[134];    
  assign wireOut[141] = wireIn[142];    
  assign wireOut[142] = wireIn[135];    
  assign wireOut[143] = wireIn[143];    
  assign wireOut[144] = wireIn[144];    
  assign wireOut[145] = wireIn[152];    
  assign wireOut[146] = wireIn[145];    
  assign wireOut[147] = wireIn[153];    
  assign wireOut[148] = wireIn[146];    
  assign wireOut[149] = wireIn[154];    
  assign wireOut[150] = wireIn[147];    
  assign wireOut[151] = wireIn[155];    
  assign wireOut[152] = wireIn[148];    
  assign wireOut[153] = wireIn[156];    
  assign wireOut[154] = wireIn[149];    
  assign wireOut[155] = wireIn[157];    
  assign wireOut[156] = wireIn[150];    
  assign wireOut[157] = wireIn[158];    
  assign wireOut[158] = wireIn[151];    
  assign wireOut[159] = wireIn[159];    
  assign wireOut[160] = wireIn[160];    
  assign wireOut[161] = wireIn[168];    
  assign wireOut[162] = wireIn[161];    
  assign wireOut[163] = wireIn[169];    
  assign wireOut[164] = wireIn[162];    
  assign wireOut[165] = wireIn[170];    
  assign wireOut[166] = wireIn[163];    
  assign wireOut[167] = wireIn[171];    
  assign wireOut[168] = wireIn[164];    
  assign wireOut[169] = wireIn[172];    
  assign wireOut[170] = wireIn[165];    
  assign wireOut[171] = wireIn[173];    
  assign wireOut[172] = wireIn[166];    
  assign wireOut[173] = wireIn[174];    
  assign wireOut[174] = wireIn[167];    
  assign wireOut[175] = wireIn[175];    
  assign wireOut[176] = wireIn[176];    
  assign wireOut[177] = wireIn[184];    
  assign wireOut[178] = wireIn[177];    
  assign wireOut[179] = wireIn[185];    
  assign wireOut[180] = wireIn[178];    
  assign wireOut[181] = wireIn[186];    
  assign wireOut[182] = wireIn[179];    
  assign wireOut[183] = wireIn[187];    
  assign wireOut[184] = wireIn[180];    
  assign wireOut[185] = wireIn[188];    
  assign wireOut[186] = wireIn[181];    
  assign wireOut[187] = wireIn[189];    
  assign wireOut[188] = wireIn[182];    
  assign wireOut[189] = wireIn[190];    
  assign wireOut[190] = wireIn[183];    
  assign wireOut[191] = wireIn[191];    
  assign wireOut[192] = wireIn[192];    
  assign wireOut[193] = wireIn[200];    
  assign wireOut[194] = wireIn[193];    
  assign wireOut[195] = wireIn[201];    
  assign wireOut[196] = wireIn[194];    
  assign wireOut[197] = wireIn[202];    
  assign wireOut[198] = wireIn[195];    
  assign wireOut[199] = wireIn[203];    
  assign wireOut[200] = wireIn[196];    
  assign wireOut[201] = wireIn[204];    
  assign wireOut[202] = wireIn[197];    
  assign wireOut[203] = wireIn[205];    
  assign wireOut[204] = wireIn[198];    
  assign wireOut[205] = wireIn[206];    
  assign wireOut[206] = wireIn[199];    
  assign wireOut[207] = wireIn[207];    
  assign wireOut[208] = wireIn[208];    
  assign wireOut[209] = wireIn[216];    
  assign wireOut[210] = wireIn[209];    
  assign wireOut[211] = wireIn[217];    
  assign wireOut[212] = wireIn[210];    
  assign wireOut[213] = wireIn[218];    
  assign wireOut[214] = wireIn[211];    
  assign wireOut[215] = wireIn[219];    
  assign wireOut[216] = wireIn[212];    
  assign wireOut[217] = wireIn[220];    
  assign wireOut[218] = wireIn[213];    
  assign wireOut[219] = wireIn[221];    
  assign wireOut[220] = wireIn[214];    
  assign wireOut[221] = wireIn[222];    
  assign wireOut[222] = wireIn[215];    
  assign wireOut[223] = wireIn[223];    
  assign wireOut[224] = wireIn[224];    
  assign wireOut[225] = wireIn[232];    
  assign wireOut[226] = wireIn[225];    
  assign wireOut[227] = wireIn[233];    
  assign wireOut[228] = wireIn[226];    
  assign wireOut[229] = wireIn[234];    
  assign wireOut[230] = wireIn[227];    
  assign wireOut[231] = wireIn[235];    
  assign wireOut[232] = wireIn[228];    
  assign wireOut[233] = wireIn[236];    
  assign wireOut[234] = wireIn[229];    
  assign wireOut[235] = wireIn[237];    
  assign wireOut[236] = wireIn[230];    
  assign wireOut[237] = wireIn[238];    
  assign wireOut[238] = wireIn[231];    
  assign wireOut[239] = wireIn[239];    
  assign wireOut[240] = wireIn[240];    
  assign wireOut[241] = wireIn[248];    
  assign wireOut[242] = wireIn[241];    
  assign wireOut[243] = wireIn[249];    
  assign wireOut[244] = wireIn[242];    
  assign wireOut[245] = wireIn[250];    
  assign wireOut[246] = wireIn[243];    
  assign wireOut[247] = wireIn[251];    
  assign wireOut[248] = wireIn[244];    
  assign wireOut[249] = wireIn[252];    
  assign wireOut[250] = wireIn[245];    
  assign wireOut[251] = wireIn[253];    
  assign wireOut[252] = wireIn[246];    
  assign wireOut[253] = wireIn[254];    
  assign wireOut[254] = wireIn[247];    
  assign wireOut[255] = wireIn[255];    
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module switches_stage_st5_0_R(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
ctrl,                            
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;                   
  input [128-1:0] ctrl;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  switch_2_2 switch_inst_0(.inData_0(wireIn[0]), .inData_1(wireIn[1]), .outData_0(wireOut[0]), .outData_1(wireOut[1]), .ctrl(ctrl[0]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_1(.inData_0(wireIn[2]), .inData_1(wireIn[3]), .outData_0(wireOut[2]), .outData_1(wireOut[3]), .ctrl(ctrl[1]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_2(.inData_0(wireIn[4]), .inData_1(wireIn[5]), .outData_0(wireOut[4]), .outData_1(wireOut[5]), .ctrl(ctrl[2]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_3(.inData_0(wireIn[6]), .inData_1(wireIn[7]), .outData_0(wireOut[6]), .outData_1(wireOut[7]), .ctrl(ctrl[3]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_4(.inData_0(wireIn[8]), .inData_1(wireIn[9]), .outData_0(wireOut[8]), .outData_1(wireOut[9]), .ctrl(ctrl[4]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_5(.inData_0(wireIn[10]), .inData_1(wireIn[11]), .outData_0(wireOut[10]), .outData_1(wireOut[11]), .ctrl(ctrl[5]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_6(.inData_0(wireIn[12]), .inData_1(wireIn[13]), .outData_0(wireOut[12]), .outData_1(wireOut[13]), .ctrl(ctrl[6]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_7(.inData_0(wireIn[14]), .inData_1(wireIn[15]), .outData_0(wireOut[14]), .outData_1(wireOut[15]), .ctrl(ctrl[7]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_8(.inData_0(wireIn[16]), .inData_1(wireIn[17]), .outData_0(wireOut[16]), .outData_1(wireOut[17]), .ctrl(ctrl[8]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_9(.inData_0(wireIn[18]), .inData_1(wireIn[19]), .outData_0(wireOut[18]), .outData_1(wireOut[19]), .ctrl(ctrl[9]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_10(.inData_0(wireIn[20]), .inData_1(wireIn[21]), .outData_0(wireOut[20]), .outData_1(wireOut[21]), .ctrl(ctrl[10]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_11(.inData_0(wireIn[22]), .inData_1(wireIn[23]), .outData_0(wireOut[22]), .outData_1(wireOut[23]), .ctrl(ctrl[11]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_12(.inData_0(wireIn[24]), .inData_1(wireIn[25]), .outData_0(wireOut[24]), .outData_1(wireOut[25]), .ctrl(ctrl[12]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_13(.inData_0(wireIn[26]), .inData_1(wireIn[27]), .outData_0(wireOut[26]), .outData_1(wireOut[27]), .ctrl(ctrl[13]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_14(.inData_0(wireIn[28]), .inData_1(wireIn[29]), .outData_0(wireOut[28]), .outData_1(wireOut[29]), .ctrl(ctrl[14]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_15(.inData_0(wireIn[30]), .inData_1(wireIn[31]), .outData_0(wireOut[30]), .outData_1(wireOut[31]), .ctrl(ctrl[15]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_16(.inData_0(wireIn[32]), .inData_1(wireIn[33]), .outData_0(wireOut[32]), .outData_1(wireOut[33]), .ctrl(ctrl[16]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_17(.inData_0(wireIn[34]), .inData_1(wireIn[35]), .outData_0(wireOut[34]), .outData_1(wireOut[35]), .ctrl(ctrl[17]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_18(.inData_0(wireIn[36]), .inData_1(wireIn[37]), .outData_0(wireOut[36]), .outData_1(wireOut[37]), .ctrl(ctrl[18]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_19(.inData_0(wireIn[38]), .inData_1(wireIn[39]), .outData_0(wireOut[38]), .outData_1(wireOut[39]), .ctrl(ctrl[19]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_20(.inData_0(wireIn[40]), .inData_1(wireIn[41]), .outData_0(wireOut[40]), .outData_1(wireOut[41]), .ctrl(ctrl[20]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_21(.inData_0(wireIn[42]), .inData_1(wireIn[43]), .outData_0(wireOut[42]), .outData_1(wireOut[43]), .ctrl(ctrl[21]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_22(.inData_0(wireIn[44]), .inData_1(wireIn[45]), .outData_0(wireOut[44]), .outData_1(wireOut[45]), .ctrl(ctrl[22]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_23(.inData_0(wireIn[46]), .inData_1(wireIn[47]), .outData_0(wireOut[46]), .outData_1(wireOut[47]), .ctrl(ctrl[23]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_24(.inData_0(wireIn[48]), .inData_1(wireIn[49]), .outData_0(wireOut[48]), .outData_1(wireOut[49]), .ctrl(ctrl[24]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_25(.inData_0(wireIn[50]), .inData_1(wireIn[51]), .outData_0(wireOut[50]), .outData_1(wireOut[51]), .ctrl(ctrl[25]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_26(.inData_0(wireIn[52]), .inData_1(wireIn[53]), .outData_0(wireOut[52]), .outData_1(wireOut[53]), .ctrl(ctrl[26]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_27(.inData_0(wireIn[54]), .inData_1(wireIn[55]), .outData_0(wireOut[54]), .outData_1(wireOut[55]), .ctrl(ctrl[27]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_28(.inData_0(wireIn[56]), .inData_1(wireIn[57]), .outData_0(wireOut[56]), .outData_1(wireOut[57]), .ctrl(ctrl[28]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_29(.inData_0(wireIn[58]), .inData_1(wireIn[59]), .outData_0(wireOut[58]), .outData_1(wireOut[59]), .ctrl(ctrl[29]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_30(.inData_0(wireIn[60]), .inData_1(wireIn[61]), .outData_0(wireOut[60]), .outData_1(wireOut[61]), .ctrl(ctrl[30]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_31(.inData_0(wireIn[62]), .inData_1(wireIn[63]), .outData_0(wireOut[62]), .outData_1(wireOut[63]), .ctrl(ctrl[31]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_32(.inData_0(wireIn[64]), .inData_1(wireIn[65]), .outData_0(wireOut[64]), .outData_1(wireOut[65]), .ctrl(ctrl[32]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_33(.inData_0(wireIn[66]), .inData_1(wireIn[67]), .outData_0(wireOut[66]), .outData_1(wireOut[67]), .ctrl(ctrl[33]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_34(.inData_0(wireIn[68]), .inData_1(wireIn[69]), .outData_0(wireOut[68]), .outData_1(wireOut[69]), .ctrl(ctrl[34]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_35(.inData_0(wireIn[70]), .inData_1(wireIn[71]), .outData_0(wireOut[70]), .outData_1(wireOut[71]), .ctrl(ctrl[35]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_36(.inData_0(wireIn[72]), .inData_1(wireIn[73]), .outData_0(wireOut[72]), .outData_1(wireOut[73]), .ctrl(ctrl[36]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_37(.inData_0(wireIn[74]), .inData_1(wireIn[75]), .outData_0(wireOut[74]), .outData_1(wireOut[75]), .ctrl(ctrl[37]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_38(.inData_0(wireIn[76]), .inData_1(wireIn[77]), .outData_0(wireOut[76]), .outData_1(wireOut[77]), .ctrl(ctrl[38]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_39(.inData_0(wireIn[78]), .inData_1(wireIn[79]), .outData_0(wireOut[78]), .outData_1(wireOut[79]), .ctrl(ctrl[39]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_40(.inData_0(wireIn[80]), .inData_1(wireIn[81]), .outData_0(wireOut[80]), .outData_1(wireOut[81]), .ctrl(ctrl[40]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_41(.inData_0(wireIn[82]), .inData_1(wireIn[83]), .outData_0(wireOut[82]), .outData_1(wireOut[83]), .ctrl(ctrl[41]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_42(.inData_0(wireIn[84]), .inData_1(wireIn[85]), .outData_0(wireOut[84]), .outData_1(wireOut[85]), .ctrl(ctrl[42]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_43(.inData_0(wireIn[86]), .inData_1(wireIn[87]), .outData_0(wireOut[86]), .outData_1(wireOut[87]), .ctrl(ctrl[43]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_44(.inData_0(wireIn[88]), .inData_1(wireIn[89]), .outData_0(wireOut[88]), .outData_1(wireOut[89]), .ctrl(ctrl[44]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_45(.inData_0(wireIn[90]), .inData_1(wireIn[91]), .outData_0(wireOut[90]), .outData_1(wireOut[91]), .ctrl(ctrl[45]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_46(.inData_0(wireIn[92]), .inData_1(wireIn[93]), .outData_0(wireOut[92]), .outData_1(wireOut[93]), .ctrl(ctrl[46]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_47(.inData_0(wireIn[94]), .inData_1(wireIn[95]), .outData_0(wireOut[94]), .outData_1(wireOut[95]), .ctrl(ctrl[47]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_48(.inData_0(wireIn[96]), .inData_1(wireIn[97]), .outData_0(wireOut[96]), .outData_1(wireOut[97]), .ctrl(ctrl[48]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_49(.inData_0(wireIn[98]), .inData_1(wireIn[99]), .outData_0(wireOut[98]), .outData_1(wireOut[99]), .ctrl(ctrl[49]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_50(.inData_0(wireIn[100]), .inData_1(wireIn[101]), .outData_0(wireOut[100]), .outData_1(wireOut[101]), .ctrl(ctrl[50]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_51(.inData_0(wireIn[102]), .inData_1(wireIn[103]), .outData_0(wireOut[102]), .outData_1(wireOut[103]), .ctrl(ctrl[51]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_52(.inData_0(wireIn[104]), .inData_1(wireIn[105]), .outData_0(wireOut[104]), .outData_1(wireOut[105]), .ctrl(ctrl[52]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_53(.inData_0(wireIn[106]), .inData_1(wireIn[107]), .outData_0(wireOut[106]), .outData_1(wireOut[107]), .ctrl(ctrl[53]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_54(.inData_0(wireIn[108]), .inData_1(wireIn[109]), .outData_0(wireOut[108]), .outData_1(wireOut[109]), .ctrl(ctrl[54]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_55(.inData_0(wireIn[110]), .inData_1(wireIn[111]), .outData_0(wireOut[110]), .outData_1(wireOut[111]), .ctrl(ctrl[55]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_56(.inData_0(wireIn[112]), .inData_1(wireIn[113]), .outData_0(wireOut[112]), .outData_1(wireOut[113]), .ctrl(ctrl[56]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_57(.inData_0(wireIn[114]), .inData_1(wireIn[115]), .outData_0(wireOut[114]), .outData_1(wireOut[115]), .ctrl(ctrl[57]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_58(.inData_0(wireIn[116]), .inData_1(wireIn[117]), .outData_0(wireOut[116]), .outData_1(wireOut[117]), .ctrl(ctrl[58]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_59(.inData_0(wireIn[118]), .inData_1(wireIn[119]), .outData_0(wireOut[118]), .outData_1(wireOut[119]), .ctrl(ctrl[59]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_60(.inData_0(wireIn[120]), .inData_1(wireIn[121]), .outData_0(wireOut[120]), .outData_1(wireOut[121]), .ctrl(ctrl[60]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_61(.inData_0(wireIn[122]), .inData_1(wireIn[123]), .outData_0(wireOut[122]), .outData_1(wireOut[123]), .ctrl(ctrl[61]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_62(.inData_0(wireIn[124]), .inData_1(wireIn[125]), .outData_0(wireOut[124]), .outData_1(wireOut[125]), .ctrl(ctrl[62]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_63(.inData_0(wireIn[126]), .inData_1(wireIn[127]), .outData_0(wireOut[126]), .outData_1(wireOut[127]), .ctrl(ctrl[63]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_64(.inData_0(wireIn[128]), .inData_1(wireIn[129]), .outData_0(wireOut[128]), .outData_1(wireOut[129]), .ctrl(ctrl[64]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_65(.inData_0(wireIn[130]), .inData_1(wireIn[131]), .outData_0(wireOut[130]), .outData_1(wireOut[131]), .ctrl(ctrl[65]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_66(.inData_0(wireIn[132]), .inData_1(wireIn[133]), .outData_0(wireOut[132]), .outData_1(wireOut[133]), .ctrl(ctrl[66]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_67(.inData_0(wireIn[134]), .inData_1(wireIn[135]), .outData_0(wireOut[134]), .outData_1(wireOut[135]), .ctrl(ctrl[67]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_68(.inData_0(wireIn[136]), .inData_1(wireIn[137]), .outData_0(wireOut[136]), .outData_1(wireOut[137]), .ctrl(ctrl[68]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_69(.inData_0(wireIn[138]), .inData_1(wireIn[139]), .outData_0(wireOut[138]), .outData_1(wireOut[139]), .ctrl(ctrl[69]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_70(.inData_0(wireIn[140]), .inData_1(wireIn[141]), .outData_0(wireOut[140]), .outData_1(wireOut[141]), .ctrl(ctrl[70]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_71(.inData_0(wireIn[142]), .inData_1(wireIn[143]), .outData_0(wireOut[142]), .outData_1(wireOut[143]), .ctrl(ctrl[71]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_72(.inData_0(wireIn[144]), .inData_1(wireIn[145]), .outData_0(wireOut[144]), .outData_1(wireOut[145]), .ctrl(ctrl[72]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_73(.inData_0(wireIn[146]), .inData_1(wireIn[147]), .outData_0(wireOut[146]), .outData_1(wireOut[147]), .ctrl(ctrl[73]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_74(.inData_0(wireIn[148]), .inData_1(wireIn[149]), .outData_0(wireOut[148]), .outData_1(wireOut[149]), .ctrl(ctrl[74]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_75(.inData_0(wireIn[150]), .inData_1(wireIn[151]), .outData_0(wireOut[150]), .outData_1(wireOut[151]), .ctrl(ctrl[75]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_76(.inData_0(wireIn[152]), .inData_1(wireIn[153]), .outData_0(wireOut[152]), .outData_1(wireOut[153]), .ctrl(ctrl[76]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_77(.inData_0(wireIn[154]), .inData_1(wireIn[155]), .outData_0(wireOut[154]), .outData_1(wireOut[155]), .ctrl(ctrl[77]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_78(.inData_0(wireIn[156]), .inData_1(wireIn[157]), .outData_0(wireOut[156]), .outData_1(wireOut[157]), .ctrl(ctrl[78]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_79(.inData_0(wireIn[158]), .inData_1(wireIn[159]), .outData_0(wireOut[158]), .outData_1(wireOut[159]), .ctrl(ctrl[79]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_80(.inData_0(wireIn[160]), .inData_1(wireIn[161]), .outData_0(wireOut[160]), .outData_1(wireOut[161]), .ctrl(ctrl[80]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_81(.inData_0(wireIn[162]), .inData_1(wireIn[163]), .outData_0(wireOut[162]), .outData_1(wireOut[163]), .ctrl(ctrl[81]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_82(.inData_0(wireIn[164]), .inData_1(wireIn[165]), .outData_0(wireOut[164]), .outData_1(wireOut[165]), .ctrl(ctrl[82]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_83(.inData_0(wireIn[166]), .inData_1(wireIn[167]), .outData_0(wireOut[166]), .outData_1(wireOut[167]), .ctrl(ctrl[83]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_84(.inData_0(wireIn[168]), .inData_1(wireIn[169]), .outData_0(wireOut[168]), .outData_1(wireOut[169]), .ctrl(ctrl[84]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_85(.inData_0(wireIn[170]), .inData_1(wireIn[171]), .outData_0(wireOut[170]), .outData_1(wireOut[171]), .ctrl(ctrl[85]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_86(.inData_0(wireIn[172]), .inData_1(wireIn[173]), .outData_0(wireOut[172]), .outData_1(wireOut[173]), .ctrl(ctrl[86]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_87(.inData_0(wireIn[174]), .inData_1(wireIn[175]), .outData_0(wireOut[174]), .outData_1(wireOut[175]), .ctrl(ctrl[87]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_88(.inData_0(wireIn[176]), .inData_1(wireIn[177]), .outData_0(wireOut[176]), .outData_1(wireOut[177]), .ctrl(ctrl[88]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_89(.inData_0(wireIn[178]), .inData_1(wireIn[179]), .outData_0(wireOut[178]), .outData_1(wireOut[179]), .ctrl(ctrl[89]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_90(.inData_0(wireIn[180]), .inData_1(wireIn[181]), .outData_0(wireOut[180]), .outData_1(wireOut[181]), .ctrl(ctrl[90]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_91(.inData_0(wireIn[182]), .inData_1(wireIn[183]), .outData_0(wireOut[182]), .outData_1(wireOut[183]), .ctrl(ctrl[91]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_92(.inData_0(wireIn[184]), .inData_1(wireIn[185]), .outData_0(wireOut[184]), .outData_1(wireOut[185]), .ctrl(ctrl[92]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_93(.inData_0(wireIn[186]), .inData_1(wireIn[187]), .outData_0(wireOut[186]), .outData_1(wireOut[187]), .ctrl(ctrl[93]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_94(.inData_0(wireIn[188]), .inData_1(wireIn[189]), .outData_0(wireOut[188]), .outData_1(wireOut[189]), .ctrl(ctrl[94]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_95(.inData_0(wireIn[190]), .inData_1(wireIn[191]), .outData_0(wireOut[190]), .outData_1(wireOut[191]), .ctrl(ctrl[95]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_96(.inData_0(wireIn[192]), .inData_1(wireIn[193]), .outData_0(wireOut[192]), .outData_1(wireOut[193]), .ctrl(ctrl[96]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_97(.inData_0(wireIn[194]), .inData_1(wireIn[195]), .outData_0(wireOut[194]), .outData_1(wireOut[195]), .ctrl(ctrl[97]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_98(.inData_0(wireIn[196]), .inData_1(wireIn[197]), .outData_0(wireOut[196]), .outData_1(wireOut[197]), .ctrl(ctrl[98]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_99(.inData_0(wireIn[198]), .inData_1(wireIn[199]), .outData_0(wireOut[198]), .outData_1(wireOut[199]), .ctrl(ctrl[99]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_100(.inData_0(wireIn[200]), .inData_1(wireIn[201]), .outData_0(wireOut[200]), .outData_1(wireOut[201]), .ctrl(ctrl[100]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_101(.inData_0(wireIn[202]), .inData_1(wireIn[203]), .outData_0(wireOut[202]), .outData_1(wireOut[203]), .ctrl(ctrl[101]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_102(.inData_0(wireIn[204]), .inData_1(wireIn[205]), .outData_0(wireOut[204]), .outData_1(wireOut[205]), .ctrl(ctrl[102]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_103(.inData_0(wireIn[206]), .inData_1(wireIn[207]), .outData_0(wireOut[206]), .outData_1(wireOut[207]), .ctrl(ctrl[103]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_104(.inData_0(wireIn[208]), .inData_1(wireIn[209]), .outData_0(wireOut[208]), .outData_1(wireOut[209]), .ctrl(ctrl[104]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_105(.inData_0(wireIn[210]), .inData_1(wireIn[211]), .outData_0(wireOut[210]), .outData_1(wireOut[211]), .ctrl(ctrl[105]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_106(.inData_0(wireIn[212]), .inData_1(wireIn[213]), .outData_0(wireOut[212]), .outData_1(wireOut[213]), .ctrl(ctrl[106]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_107(.inData_0(wireIn[214]), .inData_1(wireIn[215]), .outData_0(wireOut[214]), .outData_1(wireOut[215]), .ctrl(ctrl[107]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_108(.inData_0(wireIn[216]), .inData_1(wireIn[217]), .outData_0(wireOut[216]), .outData_1(wireOut[217]), .ctrl(ctrl[108]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_109(.inData_0(wireIn[218]), .inData_1(wireIn[219]), .outData_0(wireOut[218]), .outData_1(wireOut[219]), .ctrl(ctrl[109]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_110(.inData_0(wireIn[220]), .inData_1(wireIn[221]), .outData_0(wireOut[220]), .outData_1(wireOut[221]), .ctrl(ctrl[110]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_111(.inData_0(wireIn[222]), .inData_1(wireIn[223]), .outData_0(wireOut[222]), .outData_1(wireOut[223]), .ctrl(ctrl[111]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_112(.inData_0(wireIn[224]), .inData_1(wireIn[225]), .outData_0(wireOut[224]), .outData_1(wireOut[225]), .ctrl(ctrl[112]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_113(.inData_0(wireIn[226]), .inData_1(wireIn[227]), .outData_0(wireOut[226]), .outData_1(wireOut[227]), .ctrl(ctrl[113]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_114(.inData_0(wireIn[228]), .inData_1(wireIn[229]), .outData_0(wireOut[228]), .outData_1(wireOut[229]), .ctrl(ctrl[114]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_115(.inData_0(wireIn[230]), .inData_1(wireIn[231]), .outData_0(wireOut[230]), .outData_1(wireOut[231]), .ctrl(ctrl[115]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_116(.inData_0(wireIn[232]), .inData_1(wireIn[233]), .outData_0(wireOut[232]), .outData_1(wireOut[233]), .ctrl(ctrl[116]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_117(.inData_0(wireIn[234]), .inData_1(wireIn[235]), .outData_0(wireOut[234]), .outData_1(wireOut[235]), .ctrl(ctrl[117]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_118(.inData_0(wireIn[236]), .inData_1(wireIn[237]), .outData_0(wireOut[236]), .outData_1(wireOut[237]), .ctrl(ctrl[118]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_119(.inData_0(wireIn[238]), .inData_1(wireIn[239]), .outData_0(wireOut[238]), .outData_1(wireOut[239]), .ctrl(ctrl[119]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_120(.inData_0(wireIn[240]), .inData_1(wireIn[241]), .outData_0(wireOut[240]), .outData_1(wireOut[241]), .ctrl(ctrl[120]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_121(.inData_0(wireIn[242]), .inData_1(wireIn[243]), .outData_0(wireOut[242]), .outData_1(wireOut[243]), .ctrl(ctrl[121]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_122(.inData_0(wireIn[244]), .inData_1(wireIn[245]), .outData_0(wireOut[244]), .outData_1(wireOut[245]), .ctrl(ctrl[122]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_123(.inData_0(wireIn[246]), .inData_1(wireIn[247]), .outData_0(wireOut[246]), .outData_1(wireOut[247]), .ctrl(ctrl[123]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_124(.inData_0(wireIn[248]), .inData_1(wireIn[249]), .outData_0(wireOut[248]), .outData_1(wireOut[249]), .ctrl(ctrl[124]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_125(.inData_0(wireIn[250]), .inData_1(wireIn[251]), .outData_0(wireOut[250]), .outData_1(wireOut[251]), .ctrl(ctrl[125]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_126(.inData_0(wireIn[252]), .inData_1(wireIn[253]), .outData_0(wireOut[252]), .outData_1(wireOut[253]), .ctrl(ctrl[126]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_127(.inData_0(wireIn[254]), .inData_1(wireIn[255]), .outData_0(wireOut[254]), .outData_1(wireOut[255]), .ctrl(ctrl[127]), .clk(clk), .rst(rst));
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module wireCon_dp256_st5_R(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  assign wireOut[0] = wireIn[0];    
  assign wireOut[1] = wireIn[4];    
  assign wireOut[2] = wireIn[1];    
  assign wireOut[3] = wireIn[5];    
  assign wireOut[4] = wireIn[2];    
  assign wireOut[5] = wireIn[6];    
  assign wireOut[6] = wireIn[3];    
  assign wireOut[7] = wireIn[7];    
  assign wireOut[8] = wireIn[8];    
  assign wireOut[9] = wireIn[12];    
  assign wireOut[10] = wireIn[9];    
  assign wireOut[11] = wireIn[13];    
  assign wireOut[12] = wireIn[10];    
  assign wireOut[13] = wireIn[14];    
  assign wireOut[14] = wireIn[11];    
  assign wireOut[15] = wireIn[15];    
  assign wireOut[16] = wireIn[16];    
  assign wireOut[17] = wireIn[20];    
  assign wireOut[18] = wireIn[17];    
  assign wireOut[19] = wireIn[21];    
  assign wireOut[20] = wireIn[18];    
  assign wireOut[21] = wireIn[22];    
  assign wireOut[22] = wireIn[19];    
  assign wireOut[23] = wireIn[23];    
  assign wireOut[24] = wireIn[24];    
  assign wireOut[25] = wireIn[28];    
  assign wireOut[26] = wireIn[25];    
  assign wireOut[27] = wireIn[29];    
  assign wireOut[28] = wireIn[26];    
  assign wireOut[29] = wireIn[30];    
  assign wireOut[30] = wireIn[27];    
  assign wireOut[31] = wireIn[31];    
  assign wireOut[32] = wireIn[32];    
  assign wireOut[33] = wireIn[36];    
  assign wireOut[34] = wireIn[33];    
  assign wireOut[35] = wireIn[37];    
  assign wireOut[36] = wireIn[34];    
  assign wireOut[37] = wireIn[38];    
  assign wireOut[38] = wireIn[35];    
  assign wireOut[39] = wireIn[39];    
  assign wireOut[40] = wireIn[40];    
  assign wireOut[41] = wireIn[44];    
  assign wireOut[42] = wireIn[41];    
  assign wireOut[43] = wireIn[45];    
  assign wireOut[44] = wireIn[42];    
  assign wireOut[45] = wireIn[46];    
  assign wireOut[46] = wireIn[43];    
  assign wireOut[47] = wireIn[47];    
  assign wireOut[48] = wireIn[48];    
  assign wireOut[49] = wireIn[52];    
  assign wireOut[50] = wireIn[49];    
  assign wireOut[51] = wireIn[53];    
  assign wireOut[52] = wireIn[50];    
  assign wireOut[53] = wireIn[54];    
  assign wireOut[54] = wireIn[51];    
  assign wireOut[55] = wireIn[55];    
  assign wireOut[56] = wireIn[56];    
  assign wireOut[57] = wireIn[60];    
  assign wireOut[58] = wireIn[57];    
  assign wireOut[59] = wireIn[61];    
  assign wireOut[60] = wireIn[58];    
  assign wireOut[61] = wireIn[62];    
  assign wireOut[62] = wireIn[59];    
  assign wireOut[63] = wireIn[63];    
  assign wireOut[64] = wireIn[64];    
  assign wireOut[65] = wireIn[68];    
  assign wireOut[66] = wireIn[65];    
  assign wireOut[67] = wireIn[69];    
  assign wireOut[68] = wireIn[66];    
  assign wireOut[69] = wireIn[70];    
  assign wireOut[70] = wireIn[67];    
  assign wireOut[71] = wireIn[71];    
  assign wireOut[72] = wireIn[72];    
  assign wireOut[73] = wireIn[76];    
  assign wireOut[74] = wireIn[73];    
  assign wireOut[75] = wireIn[77];    
  assign wireOut[76] = wireIn[74];    
  assign wireOut[77] = wireIn[78];    
  assign wireOut[78] = wireIn[75];    
  assign wireOut[79] = wireIn[79];    
  assign wireOut[80] = wireIn[80];    
  assign wireOut[81] = wireIn[84];    
  assign wireOut[82] = wireIn[81];    
  assign wireOut[83] = wireIn[85];    
  assign wireOut[84] = wireIn[82];    
  assign wireOut[85] = wireIn[86];    
  assign wireOut[86] = wireIn[83];    
  assign wireOut[87] = wireIn[87];    
  assign wireOut[88] = wireIn[88];    
  assign wireOut[89] = wireIn[92];    
  assign wireOut[90] = wireIn[89];    
  assign wireOut[91] = wireIn[93];    
  assign wireOut[92] = wireIn[90];    
  assign wireOut[93] = wireIn[94];    
  assign wireOut[94] = wireIn[91];    
  assign wireOut[95] = wireIn[95];    
  assign wireOut[96] = wireIn[96];    
  assign wireOut[97] = wireIn[100];    
  assign wireOut[98] = wireIn[97];    
  assign wireOut[99] = wireIn[101];    
  assign wireOut[100] = wireIn[98];    
  assign wireOut[101] = wireIn[102];    
  assign wireOut[102] = wireIn[99];    
  assign wireOut[103] = wireIn[103];    
  assign wireOut[104] = wireIn[104];    
  assign wireOut[105] = wireIn[108];    
  assign wireOut[106] = wireIn[105];    
  assign wireOut[107] = wireIn[109];    
  assign wireOut[108] = wireIn[106];    
  assign wireOut[109] = wireIn[110];    
  assign wireOut[110] = wireIn[107];    
  assign wireOut[111] = wireIn[111];    
  assign wireOut[112] = wireIn[112];    
  assign wireOut[113] = wireIn[116];    
  assign wireOut[114] = wireIn[113];    
  assign wireOut[115] = wireIn[117];    
  assign wireOut[116] = wireIn[114];    
  assign wireOut[117] = wireIn[118];    
  assign wireOut[118] = wireIn[115];    
  assign wireOut[119] = wireIn[119];    
  assign wireOut[120] = wireIn[120];    
  assign wireOut[121] = wireIn[124];    
  assign wireOut[122] = wireIn[121];    
  assign wireOut[123] = wireIn[125];    
  assign wireOut[124] = wireIn[122];    
  assign wireOut[125] = wireIn[126];    
  assign wireOut[126] = wireIn[123];    
  assign wireOut[127] = wireIn[127];    
  assign wireOut[128] = wireIn[128];    
  assign wireOut[129] = wireIn[132];    
  assign wireOut[130] = wireIn[129];    
  assign wireOut[131] = wireIn[133];    
  assign wireOut[132] = wireIn[130];    
  assign wireOut[133] = wireIn[134];    
  assign wireOut[134] = wireIn[131];    
  assign wireOut[135] = wireIn[135];    
  assign wireOut[136] = wireIn[136];    
  assign wireOut[137] = wireIn[140];    
  assign wireOut[138] = wireIn[137];    
  assign wireOut[139] = wireIn[141];    
  assign wireOut[140] = wireIn[138];    
  assign wireOut[141] = wireIn[142];    
  assign wireOut[142] = wireIn[139];    
  assign wireOut[143] = wireIn[143];    
  assign wireOut[144] = wireIn[144];    
  assign wireOut[145] = wireIn[148];    
  assign wireOut[146] = wireIn[145];    
  assign wireOut[147] = wireIn[149];    
  assign wireOut[148] = wireIn[146];    
  assign wireOut[149] = wireIn[150];    
  assign wireOut[150] = wireIn[147];    
  assign wireOut[151] = wireIn[151];    
  assign wireOut[152] = wireIn[152];    
  assign wireOut[153] = wireIn[156];    
  assign wireOut[154] = wireIn[153];    
  assign wireOut[155] = wireIn[157];    
  assign wireOut[156] = wireIn[154];    
  assign wireOut[157] = wireIn[158];    
  assign wireOut[158] = wireIn[155];    
  assign wireOut[159] = wireIn[159];    
  assign wireOut[160] = wireIn[160];    
  assign wireOut[161] = wireIn[164];    
  assign wireOut[162] = wireIn[161];    
  assign wireOut[163] = wireIn[165];    
  assign wireOut[164] = wireIn[162];    
  assign wireOut[165] = wireIn[166];    
  assign wireOut[166] = wireIn[163];    
  assign wireOut[167] = wireIn[167];    
  assign wireOut[168] = wireIn[168];    
  assign wireOut[169] = wireIn[172];    
  assign wireOut[170] = wireIn[169];    
  assign wireOut[171] = wireIn[173];    
  assign wireOut[172] = wireIn[170];    
  assign wireOut[173] = wireIn[174];    
  assign wireOut[174] = wireIn[171];    
  assign wireOut[175] = wireIn[175];    
  assign wireOut[176] = wireIn[176];    
  assign wireOut[177] = wireIn[180];    
  assign wireOut[178] = wireIn[177];    
  assign wireOut[179] = wireIn[181];    
  assign wireOut[180] = wireIn[178];    
  assign wireOut[181] = wireIn[182];    
  assign wireOut[182] = wireIn[179];    
  assign wireOut[183] = wireIn[183];    
  assign wireOut[184] = wireIn[184];    
  assign wireOut[185] = wireIn[188];    
  assign wireOut[186] = wireIn[185];    
  assign wireOut[187] = wireIn[189];    
  assign wireOut[188] = wireIn[186];    
  assign wireOut[189] = wireIn[190];    
  assign wireOut[190] = wireIn[187];    
  assign wireOut[191] = wireIn[191];    
  assign wireOut[192] = wireIn[192];    
  assign wireOut[193] = wireIn[196];    
  assign wireOut[194] = wireIn[193];    
  assign wireOut[195] = wireIn[197];    
  assign wireOut[196] = wireIn[194];    
  assign wireOut[197] = wireIn[198];    
  assign wireOut[198] = wireIn[195];    
  assign wireOut[199] = wireIn[199];    
  assign wireOut[200] = wireIn[200];    
  assign wireOut[201] = wireIn[204];    
  assign wireOut[202] = wireIn[201];    
  assign wireOut[203] = wireIn[205];    
  assign wireOut[204] = wireIn[202];    
  assign wireOut[205] = wireIn[206];    
  assign wireOut[206] = wireIn[203];    
  assign wireOut[207] = wireIn[207];    
  assign wireOut[208] = wireIn[208];    
  assign wireOut[209] = wireIn[212];    
  assign wireOut[210] = wireIn[209];    
  assign wireOut[211] = wireIn[213];    
  assign wireOut[212] = wireIn[210];    
  assign wireOut[213] = wireIn[214];    
  assign wireOut[214] = wireIn[211];    
  assign wireOut[215] = wireIn[215];    
  assign wireOut[216] = wireIn[216];    
  assign wireOut[217] = wireIn[220];    
  assign wireOut[218] = wireIn[217];    
  assign wireOut[219] = wireIn[221];    
  assign wireOut[220] = wireIn[218];    
  assign wireOut[221] = wireIn[222];    
  assign wireOut[222] = wireIn[219];    
  assign wireOut[223] = wireIn[223];    
  assign wireOut[224] = wireIn[224];    
  assign wireOut[225] = wireIn[228];    
  assign wireOut[226] = wireIn[225];    
  assign wireOut[227] = wireIn[229];    
  assign wireOut[228] = wireIn[226];    
  assign wireOut[229] = wireIn[230];    
  assign wireOut[230] = wireIn[227];    
  assign wireOut[231] = wireIn[231];    
  assign wireOut[232] = wireIn[232];    
  assign wireOut[233] = wireIn[236];    
  assign wireOut[234] = wireIn[233];    
  assign wireOut[235] = wireIn[237];    
  assign wireOut[236] = wireIn[234];    
  assign wireOut[237] = wireIn[238];    
  assign wireOut[238] = wireIn[235];    
  assign wireOut[239] = wireIn[239];    
  assign wireOut[240] = wireIn[240];    
  assign wireOut[241] = wireIn[244];    
  assign wireOut[242] = wireIn[241];    
  assign wireOut[243] = wireIn[245];    
  assign wireOut[244] = wireIn[242];    
  assign wireOut[245] = wireIn[246];    
  assign wireOut[246] = wireIn[243];    
  assign wireOut[247] = wireIn[247];    
  assign wireOut[248] = wireIn[248];    
  assign wireOut[249] = wireIn[252];    
  assign wireOut[250] = wireIn[249];    
  assign wireOut[251] = wireIn[253];    
  assign wireOut[252] = wireIn[250];    
  assign wireOut[253] = wireIn[254];    
  assign wireOut[254] = wireIn[251];    
  assign wireOut[255] = wireIn[255];    
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module switches_stage_st6_0_R(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
ctrl,                            
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;                   
  input [128-1:0] ctrl;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  switch_2_2 switch_inst_0(.inData_0(wireIn[0]), .inData_1(wireIn[1]), .outData_0(wireOut[0]), .outData_1(wireOut[1]), .ctrl(ctrl[0]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_1(.inData_0(wireIn[2]), .inData_1(wireIn[3]), .outData_0(wireOut[2]), .outData_1(wireOut[3]), .ctrl(ctrl[1]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_2(.inData_0(wireIn[4]), .inData_1(wireIn[5]), .outData_0(wireOut[4]), .outData_1(wireOut[5]), .ctrl(ctrl[2]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_3(.inData_0(wireIn[6]), .inData_1(wireIn[7]), .outData_0(wireOut[6]), .outData_1(wireOut[7]), .ctrl(ctrl[3]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_4(.inData_0(wireIn[8]), .inData_1(wireIn[9]), .outData_0(wireOut[8]), .outData_1(wireOut[9]), .ctrl(ctrl[4]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_5(.inData_0(wireIn[10]), .inData_1(wireIn[11]), .outData_0(wireOut[10]), .outData_1(wireOut[11]), .ctrl(ctrl[5]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_6(.inData_0(wireIn[12]), .inData_1(wireIn[13]), .outData_0(wireOut[12]), .outData_1(wireOut[13]), .ctrl(ctrl[6]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_7(.inData_0(wireIn[14]), .inData_1(wireIn[15]), .outData_0(wireOut[14]), .outData_1(wireOut[15]), .ctrl(ctrl[7]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_8(.inData_0(wireIn[16]), .inData_1(wireIn[17]), .outData_0(wireOut[16]), .outData_1(wireOut[17]), .ctrl(ctrl[8]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_9(.inData_0(wireIn[18]), .inData_1(wireIn[19]), .outData_0(wireOut[18]), .outData_1(wireOut[19]), .ctrl(ctrl[9]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_10(.inData_0(wireIn[20]), .inData_1(wireIn[21]), .outData_0(wireOut[20]), .outData_1(wireOut[21]), .ctrl(ctrl[10]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_11(.inData_0(wireIn[22]), .inData_1(wireIn[23]), .outData_0(wireOut[22]), .outData_1(wireOut[23]), .ctrl(ctrl[11]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_12(.inData_0(wireIn[24]), .inData_1(wireIn[25]), .outData_0(wireOut[24]), .outData_1(wireOut[25]), .ctrl(ctrl[12]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_13(.inData_0(wireIn[26]), .inData_1(wireIn[27]), .outData_0(wireOut[26]), .outData_1(wireOut[27]), .ctrl(ctrl[13]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_14(.inData_0(wireIn[28]), .inData_1(wireIn[29]), .outData_0(wireOut[28]), .outData_1(wireOut[29]), .ctrl(ctrl[14]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_15(.inData_0(wireIn[30]), .inData_1(wireIn[31]), .outData_0(wireOut[30]), .outData_1(wireOut[31]), .ctrl(ctrl[15]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_16(.inData_0(wireIn[32]), .inData_1(wireIn[33]), .outData_0(wireOut[32]), .outData_1(wireOut[33]), .ctrl(ctrl[16]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_17(.inData_0(wireIn[34]), .inData_1(wireIn[35]), .outData_0(wireOut[34]), .outData_1(wireOut[35]), .ctrl(ctrl[17]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_18(.inData_0(wireIn[36]), .inData_1(wireIn[37]), .outData_0(wireOut[36]), .outData_1(wireOut[37]), .ctrl(ctrl[18]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_19(.inData_0(wireIn[38]), .inData_1(wireIn[39]), .outData_0(wireOut[38]), .outData_1(wireOut[39]), .ctrl(ctrl[19]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_20(.inData_0(wireIn[40]), .inData_1(wireIn[41]), .outData_0(wireOut[40]), .outData_1(wireOut[41]), .ctrl(ctrl[20]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_21(.inData_0(wireIn[42]), .inData_1(wireIn[43]), .outData_0(wireOut[42]), .outData_1(wireOut[43]), .ctrl(ctrl[21]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_22(.inData_0(wireIn[44]), .inData_1(wireIn[45]), .outData_0(wireOut[44]), .outData_1(wireOut[45]), .ctrl(ctrl[22]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_23(.inData_0(wireIn[46]), .inData_1(wireIn[47]), .outData_0(wireOut[46]), .outData_1(wireOut[47]), .ctrl(ctrl[23]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_24(.inData_0(wireIn[48]), .inData_1(wireIn[49]), .outData_0(wireOut[48]), .outData_1(wireOut[49]), .ctrl(ctrl[24]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_25(.inData_0(wireIn[50]), .inData_1(wireIn[51]), .outData_0(wireOut[50]), .outData_1(wireOut[51]), .ctrl(ctrl[25]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_26(.inData_0(wireIn[52]), .inData_1(wireIn[53]), .outData_0(wireOut[52]), .outData_1(wireOut[53]), .ctrl(ctrl[26]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_27(.inData_0(wireIn[54]), .inData_1(wireIn[55]), .outData_0(wireOut[54]), .outData_1(wireOut[55]), .ctrl(ctrl[27]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_28(.inData_0(wireIn[56]), .inData_1(wireIn[57]), .outData_0(wireOut[56]), .outData_1(wireOut[57]), .ctrl(ctrl[28]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_29(.inData_0(wireIn[58]), .inData_1(wireIn[59]), .outData_0(wireOut[58]), .outData_1(wireOut[59]), .ctrl(ctrl[29]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_30(.inData_0(wireIn[60]), .inData_1(wireIn[61]), .outData_0(wireOut[60]), .outData_1(wireOut[61]), .ctrl(ctrl[30]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_31(.inData_0(wireIn[62]), .inData_1(wireIn[63]), .outData_0(wireOut[62]), .outData_1(wireOut[63]), .ctrl(ctrl[31]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_32(.inData_0(wireIn[64]), .inData_1(wireIn[65]), .outData_0(wireOut[64]), .outData_1(wireOut[65]), .ctrl(ctrl[32]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_33(.inData_0(wireIn[66]), .inData_1(wireIn[67]), .outData_0(wireOut[66]), .outData_1(wireOut[67]), .ctrl(ctrl[33]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_34(.inData_0(wireIn[68]), .inData_1(wireIn[69]), .outData_0(wireOut[68]), .outData_1(wireOut[69]), .ctrl(ctrl[34]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_35(.inData_0(wireIn[70]), .inData_1(wireIn[71]), .outData_0(wireOut[70]), .outData_1(wireOut[71]), .ctrl(ctrl[35]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_36(.inData_0(wireIn[72]), .inData_1(wireIn[73]), .outData_0(wireOut[72]), .outData_1(wireOut[73]), .ctrl(ctrl[36]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_37(.inData_0(wireIn[74]), .inData_1(wireIn[75]), .outData_0(wireOut[74]), .outData_1(wireOut[75]), .ctrl(ctrl[37]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_38(.inData_0(wireIn[76]), .inData_1(wireIn[77]), .outData_0(wireOut[76]), .outData_1(wireOut[77]), .ctrl(ctrl[38]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_39(.inData_0(wireIn[78]), .inData_1(wireIn[79]), .outData_0(wireOut[78]), .outData_1(wireOut[79]), .ctrl(ctrl[39]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_40(.inData_0(wireIn[80]), .inData_1(wireIn[81]), .outData_0(wireOut[80]), .outData_1(wireOut[81]), .ctrl(ctrl[40]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_41(.inData_0(wireIn[82]), .inData_1(wireIn[83]), .outData_0(wireOut[82]), .outData_1(wireOut[83]), .ctrl(ctrl[41]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_42(.inData_0(wireIn[84]), .inData_1(wireIn[85]), .outData_0(wireOut[84]), .outData_1(wireOut[85]), .ctrl(ctrl[42]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_43(.inData_0(wireIn[86]), .inData_1(wireIn[87]), .outData_0(wireOut[86]), .outData_1(wireOut[87]), .ctrl(ctrl[43]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_44(.inData_0(wireIn[88]), .inData_1(wireIn[89]), .outData_0(wireOut[88]), .outData_1(wireOut[89]), .ctrl(ctrl[44]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_45(.inData_0(wireIn[90]), .inData_1(wireIn[91]), .outData_0(wireOut[90]), .outData_1(wireOut[91]), .ctrl(ctrl[45]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_46(.inData_0(wireIn[92]), .inData_1(wireIn[93]), .outData_0(wireOut[92]), .outData_1(wireOut[93]), .ctrl(ctrl[46]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_47(.inData_0(wireIn[94]), .inData_1(wireIn[95]), .outData_0(wireOut[94]), .outData_1(wireOut[95]), .ctrl(ctrl[47]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_48(.inData_0(wireIn[96]), .inData_1(wireIn[97]), .outData_0(wireOut[96]), .outData_1(wireOut[97]), .ctrl(ctrl[48]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_49(.inData_0(wireIn[98]), .inData_1(wireIn[99]), .outData_0(wireOut[98]), .outData_1(wireOut[99]), .ctrl(ctrl[49]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_50(.inData_0(wireIn[100]), .inData_1(wireIn[101]), .outData_0(wireOut[100]), .outData_1(wireOut[101]), .ctrl(ctrl[50]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_51(.inData_0(wireIn[102]), .inData_1(wireIn[103]), .outData_0(wireOut[102]), .outData_1(wireOut[103]), .ctrl(ctrl[51]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_52(.inData_0(wireIn[104]), .inData_1(wireIn[105]), .outData_0(wireOut[104]), .outData_1(wireOut[105]), .ctrl(ctrl[52]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_53(.inData_0(wireIn[106]), .inData_1(wireIn[107]), .outData_0(wireOut[106]), .outData_1(wireOut[107]), .ctrl(ctrl[53]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_54(.inData_0(wireIn[108]), .inData_1(wireIn[109]), .outData_0(wireOut[108]), .outData_1(wireOut[109]), .ctrl(ctrl[54]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_55(.inData_0(wireIn[110]), .inData_1(wireIn[111]), .outData_0(wireOut[110]), .outData_1(wireOut[111]), .ctrl(ctrl[55]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_56(.inData_0(wireIn[112]), .inData_1(wireIn[113]), .outData_0(wireOut[112]), .outData_1(wireOut[113]), .ctrl(ctrl[56]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_57(.inData_0(wireIn[114]), .inData_1(wireIn[115]), .outData_0(wireOut[114]), .outData_1(wireOut[115]), .ctrl(ctrl[57]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_58(.inData_0(wireIn[116]), .inData_1(wireIn[117]), .outData_0(wireOut[116]), .outData_1(wireOut[117]), .ctrl(ctrl[58]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_59(.inData_0(wireIn[118]), .inData_1(wireIn[119]), .outData_0(wireOut[118]), .outData_1(wireOut[119]), .ctrl(ctrl[59]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_60(.inData_0(wireIn[120]), .inData_1(wireIn[121]), .outData_0(wireOut[120]), .outData_1(wireOut[121]), .ctrl(ctrl[60]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_61(.inData_0(wireIn[122]), .inData_1(wireIn[123]), .outData_0(wireOut[122]), .outData_1(wireOut[123]), .ctrl(ctrl[61]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_62(.inData_0(wireIn[124]), .inData_1(wireIn[125]), .outData_0(wireOut[124]), .outData_1(wireOut[125]), .ctrl(ctrl[62]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_63(.inData_0(wireIn[126]), .inData_1(wireIn[127]), .outData_0(wireOut[126]), .outData_1(wireOut[127]), .ctrl(ctrl[63]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_64(.inData_0(wireIn[128]), .inData_1(wireIn[129]), .outData_0(wireOut[128]), .outData_1(wireOut[129]), .ctrl(ctrl[64]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_65(.inData_0(wireIn[130]), .inData_1(wireIn[131]), .outData_0(wireOut[130]), .outData_1(wireOut[131]), .ctrl(ctrl[65]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_66(.inData_0(wireIn[132]), .inData_1(wireIn[133]), .outData_0(wireOut[132]), .outData_1(wireOut[133]), .ctrl(ctrl[66]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_67(.inData_0(wireIn[134]), .inData_1(wireIn[135]), .outData_0(wireOut[134]), .outData_1(wireOut[135]), .ctrl(ctrl[67]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_68(.inData_0(wireIn[136]), .inData_1(wireIn[137]), .outData_0(wireOut[136]), .outData_1(wireOut[137]), .ctrl(ctrl[68]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_69(.inData_0(wireIn[138]), .inData_1(wireIn[139]), .outData_0(wireOut[138]), .outData_1(wireOut[139]), .ctrl(ctrl[69]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_70(.inData_0(wireIn[140]), .inData_1(wireIn[141]), .outData_0(wireOut[140]), .outData_1(wireOut[141]), .ctrl(ctrl[70]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_71(.inData_0(wireIn[142]), .inData_1(wireIn[143]), .outData_0(wireOut[142]), .outData_1(wireOut[143]), .ctrl(ctrl[71]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_72(.inData_0(wireIn[144]), .inData_1(wireIn[145]), .outData_0(wireOut[144]), .outData_1(wireOut[145]), .ctrl(ctrl[72]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_73(.inData_0(wireIn[146]), .inData_1(wireIn[147]), .outData_0(wireOut[146]), .outData_1(wireOut[147]), .ctrl(ctrl[73]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_74(.inData_0(wireIn[148]), .inData_1(wireIn[149]), .outData_0(wireOut[148]), .outData_1(wireOut[149]), .ctrl(ctrl[74]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_75(.inData_0(wireIn[150]), .inData_1(wireIn[151]), .outData_0(wireOut[150]), .outData_1(wireOut[151]), .ctrl(ctrl[75]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_76(.inData_0(wireIn[152]), .inData_1(wireIn[153]), .outData_0(wireOut[152]), .outData_1(wireOut[153]), .ctrl(ctrl[76]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_77(.inData_0(wireIn[154]), .inData_1(wireIn[155]), .outData_0(wireOut[154]), .outData_1(wireOut[155]), .ctrl(ctrl[77]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_78(.inData_0(wireIn[156]), .inData_1(wireIn[157]), .outData_0(wireOut[156]), .outData_1(wireOut[157]), .ctrl(ctrl[78]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_79(.inData_0(wireIn[158]), .inData_1(wireIn[159]), .outData_0(wireOut[158]), .outData_1(wireOut[159]), .ctrl(ctrl[79]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_80(.inData_0(wireIn[160]), .inData_1(wireIn[161]), .outData_0(wireOut[160]), .outData_1(wireOut[161]), .ctrl(ctrl[80]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_81(.inData_0(wireIn[162]), .inData_1(wireIn[163]), .outData_0(wireOut[162]), .outData_1(wireOut[163]), .ctrl(ctrl[81]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_82(.inData_0(wireIn[164]), .inData_1(wireIn[165]), .outData_0(wireOut[164]), .outData_1(wireOut[165]), .ctrl(ctrl[82]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_83(.inData_0(wireIn[166]), .inData_1(wireIn[167]), .outData_0(wireOut[166]), .outData_1(wireOut[167]), .ctrl(ctrl[83]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_84(.inData_0(wireIn[168]), .inData_1(wireIn[169]), .outData_0(wireOut[168]), .outData_1(wireOut[169]), .ctrl(ctrl[84]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_85(.inData_0(wireIn[170]), .inData_1(wireIn[171]), .outData_0(wireOut[170]), .outData_1(wireOut[171]), .ctrl(ctrl[85]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_86(.inData_0(wireIn[172]), .inData_1(wireIn[173]), .outData_0(wireOut[172]), .outData_1(wireOut[173]), .ctrl(ctrl[86]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_87(.inData_0(wireIn[174]), .inData_1(wireIn[175]), .outData_0(wireOut[174]), .outData_1(wireOut[175]), .ctrl(ctrl[87]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_88(.inData_0(wireIn[176]), .inData_1(wireIn[177]), .outData_0(wireOut[176]), .outData_1(wireOut[177]), .ctrl(ctrl[88]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_89(.inData_0(wireIn[178]), .inData_1(wireIn[179]), .outData_0(wireOut[178]), .outData_1(wireOut[179]), .ctrl(ctrl[89]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_90(.inData_0(wireIn[180]), .inData_1(wireIn[181]), .outData_0(wireOut[180]), .outData_1(wireOut[181]), .ctrl(ctrl[90]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_91(.inData_0(wireIn[182]), .inData_1(wireIn[183]), .outData_0(wireOut[182]), .outData_1(wireOut[183]), .ctrl(ctrl[91]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_92(.inData_0(wireIn[184]), .inData_1(wireIn[185]), .outData_0(wireOut[184]), .outData_1(wireOut[185]), .ctrl(ctrl[92]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_93(.inData_0(wireIn[186]), .inData_1(wireIn[187]), .outData_0(wireOut[186]), .outData_1(wireOut[187]), .ctrl(ctrl[93]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_94(.inData_0(wireIn[188]), .inData_1(wireIn[189]), .outData_0(wireOut[188]), .outData_1(wireOut[189]), .ctrl(ctrl[94]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_95(.inData_0(wireIn[190]), .inData_1(wireIn[191]), .outData_0(wireOut[190]), .outData_1(wireOut[191]), .ctrl(ctrl[95]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_96(.inData_0(wireIn[192]), .inData_1(wireIn[193]), .outData_0(wireOut[192]), .outData_1(wireOut[193]), .ctrl(ctrl[96]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_97(.inData_0(wireIn[194]), .inData_1(wireIn[195]), .outData_0(wireOut[194]), .outData_1(wireOut[195]), .ctrl(ctrl[97]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_98(.inData_0(wireIn[196]), .inData_1(wireIn[197]), .outData_0(wireOut[196]), .outData_1(wireOut[197]), .ctrl(ctrl[98]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_99(.inData_0(wireIn[198]), .inData_1(wireIn[199]), .outData_0(wireOut[198]), .outData_1(wireOut[199]), .ctrl(ctrl[99]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_100(.inData_0(wireIn[200]), .inData_1(wireIn[201]), .outData_0(wireOut[200]), .outData_1(wireOut[201]), .ctrl(ctrl[100]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_101(.inData_0(wireIn[202]), .inData_1(wireIn[203]), .outData_0(wireOut[202]), .outData_1(wireOut[203]), .ctrl(ctrl[101]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_102(.inData_0(wireIn[204]), .inData_1(wireIn[205]), .outData_0(wireOut[204]), .outData_1(wireOut[205]), .ctrl(ctrl[102]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_103(.inData_0(wireIn[206]), .inData_1(wireIn[207]), .outData_0(wireOut[206]), .outData_1(wireOut[207]), .ctrl(ctrl[103]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_104(.inData_0(wireIn[208]), .inData_1(wireIn[209]), .outData_0(wireOut[208]), .outData_1(wireOut[209]), .ctrl(ctrl[104]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_105(.inData_0(wireIn[210]), .inData_1(wireIn[211]), .outData_0(wireOut[210]), .outData_1(wireOut[211]), .ctrl(ctrl[105]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_106(.inData_0(wireIn[212]), .inData_1(wireIn[213]), .outData_0(wireOut[212]), .outData_1(wireOut[213]), .ctrl(ctrl[106]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_107(.inData_0(wireIn[214]), .inData_1(wireIn[215]), .outData_0(wireOut[214]), .outData_1(wireOut[215]), .ctrl(ctrl[107]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_108(.inData_0(wireIn[216]), .inData_1(wireIn[217]), .outData_0(wireOut[216]), .outData_1(wireOut[217]), .ctrl(ctrl[108]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_109(.inData_0(wireIn[218]), .inData_1(wireIn[219]), .outData_0(wireOut[218]), .outData_1(wireOut[219]), .ctrl(ctrl[109]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_110(.inData_0(wireIn[220]), .inData_1(wireIn[221]), .outData_0(wireOut[220]), .outData_1(wireOut[221]), .ctrl(ctrl[110]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_111(.inData_0(wireIn[222]), .inData_1(wireIn[223]), .outData_0(wireOut[222]), .outData_1(wireOut[223]), .ctrl(ctrl[111]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_112(.inData_0(wireIn[224]), .inData_1(wireIn[225]), .outData_0(wireOut[224]), .outData_1(wireOut[225]), .ctrl(ctrl[112]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_113(.inData_0(wireIn[226]), .inData_1(wireIn[227]), .outData_0(wireOut[226]), .outData_1(wireOut[227]), .ctrl(ctrl[113]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_114(.inData_0(wireIn[228]), .inData_1(wireIn[229]), .outData_0(wireOut[228]), .outData_1(wireOut[229]), .ctrl(ctrl[114]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_115(.inData_0(wireIn[230]), .inData_1(wireIn[231]), .outData_0(wireOut[230]), .outData_1(wireOut[231]), .ctrl(ctrl[115]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_116(.inData_0(wireIn[232]), .inData_1(wireIn[233]), .outData_0(wireOut[232]), .outData_1(wireOut[233]), .ctrl(ctrl[116]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_117(.inData_0(wireIn[234]), .inData_1(wireIn[235]), .outData_0(wireOut[234]), .outData_1(wireOut[235]), .ctrl(ctrl[117]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_118(.inData_0(wireIn[236]), .inData_1(wireIn[237]), .outData_0(wireOut[236]), .outData_1(wireOut[237]), .ctrl(ctrl[118]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_119(.inData_0(wireIn[238]), .inData_1(wireIn[239]), .outData_0(wireOut[238]), .outData_1(wireOut[239]), .ctrl(ctrl[119]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_120(.inData_0(wireIn[240]), .inData_1(wireIn[241]), .outData_0(wireOut[240]), .outData_1(wireOut[241]), .ctrl(ctrl[120]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_121(.inData_0(wireIn[242]), .inData_1(wireIn[243]), .outData_0(wireOut[242]), .outData_1(wireOut[243]), .ctrl(ctrl[121]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_122(.inData_0(wireIn[244]), .inData_1(wireIn[245]), .outData_0(wireOut[244]), .outData_1(wireOut[245]), .ctrl(ctrl[122]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_123(.inData_0(wireIn[246]), .inData_1(wireIn[247]), .outData_0(wireOut[246]), .outData_1(wireOut[247]), .ctrl(ctrl[123]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_124(.inData_0(wireIn[248]), .inData_1(wireIn[249]), .outData_0(wireOut[248]), .outData_1(wireOut[249]), .ctrl(ctrl[124]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_125(.inData_0(wireIn[250]), .inData_1(wireIn[251]), .outData_0(wireOut[250]), .outData_1(wireOut[251]), .ctrl(ctrl[125]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_126(.inData_0(wireIn[252]), .inData_1(wireIn[253]), .outData_0(wireOut[252]), .outData_1(wireOut[253]), .ctrl(ctrl[126]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_127(.inData_0(wireIn[254]), .inData_1(wireIn[255]), .outData_0(wireOut[254]), .outData_1(wireOut[255]), .ctrl(ctrl[127]), .clk(clk), .rst(rst));
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module wireCon_dp256_st6_R(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  assign wireOut[0] = wireIn[0];    
  assign wireOut[1] = wireIn[2];    
  assign wireOut[2] = wireIn[1];    
  assign wireOut[3] = wireIn[3];    
  assign wireOut[4] = wireIn[4];    
  assign wireOut[5] = wireIn[6];    
  assign wireOut[6] = wireIn[5];    
  assign wireOut[7] = wireIn[7];    
  assign wireOut[8] = wireIn[8];    
  assign wireOut[9] = wireIn[10];    
  assign wireOut[10] = wireIn[9];    
  assign wireOut[11] = wireIn[11];    
  assign wireOut[12] = wireIn[12];    
  assign wireOut[13] = wireIn[14];    
  assign wireOut[14] = wireIn[13];    
  assign wireOut[15] = wireIn[15];    
  assign wireOut[16] = wireIn[16];    
  assign wireOut[17] = wireIn[18];    
  assign wireOut[18] = wireIn[17];    
  assign wireOut[19] = wireIn[19];    
  assign wireOut[20] = wireIn[20];    
  assign wireOut[21] = wireIn[22];    
  assign wireOut[22] = wireIn[21];    
  assign wireOut[23] = wireIn[23];    
  assign wireOut[24] = wireIn[24];    
  assign wireOut[25] = wireIn[26];    
  assign wireOut[26] = wireIn[25];    
  assign wireOut[27] = wireIn[27];    
  assign wireOut[28] = wireIn[28];    
  assign wireOut[29] = wireIn[30];    
  assign wireOut[30] = wireIn[29];    
  assign wireOut[31] = wireIn[31];    
  assign wireOut[32] = wireIn[32];    
  assign wireOut[33] = wireIn[34];    
  assign wireOut[34] = wireIn[33];    
  assign wireOut[35] = wireIn[35];    
  assign wireOut[36] = wireIn[36];    
  assign wireOut[37] = wireIn[38];    
  assign wireOut[38] = wireIn[37];    
  assign wireOut[39] = wireIn[39];    
  assign wireOut[40] = wireIn[40];    
  assign wireOut[41] = wireIn[42];    
  assign wireOut[42] = wireIn[41];    
  assign wireOut[43] = wireIn[43];    
  assign wireOut[44] = wireIn[44];    
  assign wireOut[45] = wireIn[46];    
  assign wireOut[46] = wireIn[45];    
  assign wireOut[47] = wireIn[47];    
  assign wireOut[48] = wireIn[48];    
  assign wireOut[49] = wireIn[50];    
  assign wireOut[50] = wireIn[49];    
  assign wireOut[51] = wireIn[51];    
  assign wireOut[52] = wireIn[52];    
  assign wireOut[53] = wireIn[54];    
  assign wireOut[54] = wireIn[53];    
  assign wireOut[55] = wireIn[55];    
  assign wireOut[56] = wireIn[56];    
  assign wireOut[57] = wireIn[58];    
  assign wireOut[58] = wireIn[57];    
  assign wireOut[59] = wireIn[59];    
  assign wireOut[60] = wireIn[60];    
  assign wireOut[61] = wireIn[62];    
  assign wireOut[62] = wireIn[61];    
  assign wireOut[63] = wireIn[63];    
  assign wireOut[64] = wireIn[64];    
  assign wireOut[65] = wireIn[66];    
  assign wireOut[66] = wireIn[65];    
  assign wireOut[67] = wireIn[67];    
  assign wireOut[68] = wireIn[68];    
  assign wireOut[69] = wireIn[70];    
  assign wireOut[70] = wireIn[69];    
  assign wireOut[71] = wireIn[71];    
  assign wireOut[72] = wireIn[72];    
  assign wireOut[73] = wireIn[74];    
  assign wireOut[74] = wireIn[73];    
  assign wireOut[75] = wireIn[75];    
  assign wireOut[76] = wireIn[76];    
  assign wireOut[77] = wireIn[78];    
  assign wireOut[78] = wireIn[77];    
  assign wireOut[79] = wireIn[79];    
  assign wireOut[80] = wireIn[80];    
  assign wireOut[81] = wireIn[82];    
  assign wireOut[82] = wireIn[81];    
  assign wireOut[83] = wireIn[83];    
  assign wireOut[84] = wireIn[84];    
  assign wireOut[85] = wireIn[86];    
  assign wireOut[86] = wireIn[85];    
  assign wireOut[87] = wireIn[87];    
  assign wireOut[88] = wireIn[88];    
  assign wireOut[89] = wireIn[90];    
  assign wireOut[90] = wireIn[89];    
  assign wireOut[91] = wireIn[91];    
  assign wireOut[92] = wireIn[92];    
  assign wireOut[93] = wireIn[94];    
  assign wireOut[94] = wireIn[93];    
  assign wireOut[95] = wireIn[95];    
  assign wireOut[96] = wireIn[96];    
  assign wireOut[97] = wireIn[98];    
  assign wireOut[98] = wireIn[97];    
  assign wireOut[99] = wireIn[99];    
  assign wireOut[100] = wireIn[100];    
  assign wireOut[101] = wireIn[102];    
  assign wireOut[102] = wireIn[101];    
  assign wireOut[103] = wireIn[103];    
  assign wireOut[104] = wireIn[104];    
  assign wireOut[105] = wireIn[106];    
  assign wireOut[106] = wireIn[105];    
  assign wireOut[107] = wireIn[107];    
  assign wireOut[108] = wireIn[108];    
  assign wireOut[109] = wireIn[110];    
  assign wireOut[110] = wireIn[109];    
  assign wireOut[111] = wireIn[111];    
  assign wireOut[112] = wireIn[112];    
  assign wireOut[113] = wireIn[114];    
  assign wireOut[114] = wireIn[113];    
  assign wireOut[115] = wireIn[115];    
  assign wireOut[116] = wireIn[116];    
  assign wireOut[117] = wireIn[118];    
  assign wireOut[118] = wireIn[117];    
  assign wireOut[119] = wireIn[119];    
  assign wireOut[120] = wireIn[120];    
  assign wireOut[121] = wireIn[122];    
  assign wireOut[122] = wireIn[121];    
  assign wireOut[123] = wireIn[123];    
  assign wireOut[124] = wireIn[124];    
  assign wireOut[125] = wireIn[126];    
  assign wireOut[126] = wireIn[125];    
  assign wireOut[127] = wireIn[127];    
  assign wireOut[128] = wireIn[128];    
  assign wireOut[129] = wireIn[130];    
  assign wireOut[130] = wireIn[129];    
  assign wireOut[131] = wireIn[131];    
  assign wireOut[132] = wireIn[132];    
  assign wireOut[133] = wireIn[134];    
  assign wireOut[134] = wireIn[133];    
  assign wireOut[135] = wireIn[135];    
  assign wireOut[136] = wireIn[136];    
  assign wireOut[137] = wireIn[138];    
  assign wireOut[138] = wireIn[137];    
  assign wireOut[139] = wireIn[139];    
  assign wireOut[140] = wireIn[140];    
  assign wireOut[141] = wireIn[142];    
  assign wireOut[142] = wireIn[141];    
  assign wireOut[143] = wireIn[143];    
  assign wireOut[144] = wireIn[144];    
  assign wireOut[145] = wireIn[146];    
  assign wireOut[146] = wireIn[145];    
  assign wireOut[147] = wireIn[147];    
  assign wireOut[148] = wireIn[148];    
  assign wireOut[149] = wireIn[150];    
  assign wireOut[150] = wireIn[149];    
  assign wireOut[151] = wireIn[151];    
  assign wireOut[152] = wireIn[152];    
  assign wireOut[153] = wireIn[154];    
  assign wireOut[154] = wireIn[153];    
  assign wireOut[155] = wireIn[155];    
  assign wireOut[156] = wireIn[156];    
  assign wireOut[157] = wireIn[158];    
  assign wireOut[158] = wireIn[157];    
  assign wireOut[159] = wireIn[159];    
  assign wireOut[160] = wireIn[160];    
  assign wireOut[161] = wireIn[162];    
  assign wireOut[162] = wireIn[161];    
  assign wireOut[163] = wireIn[163];    
  assign wireOut[164] = wireIn[164];    
  assign wireOut[165] = wireIn[166];    
  assign wireOut[166] = wireIn[165];    
  assign wireOut[167] = wireIn[167];    
  assign wireOut[168] = wireIn[168];    
  assign wireOut[169] = wireIn[170];    
  assign wireOut[170] = wireIn[169];    
  assign wireOut[171] = wireIn[171];    
  assign wireOut[172] = wireIn[172];    
  assign wireOut[173] = wireIn[174];    
  assign wireOut[174] = wireIn[173];    
  assign wireOut[175] = wireIn[175];    
  assign wireOut[176] = wireIn[176];    
  assign wireOut[177] = wireIn[178];    
  assign wireOut[178] = wireIn[177];    
  assign wireOut[179] = wireIn[179];    
  assign wireOut[180] = wireIn[180];    
  assign wireOut[181] = wireIn[182];    
  assign wireOut[182] = wireIn[181];    
  assign wireOut[183] = wireIn[183];    
  assign wireOut[184] = wireIn[184];    
  assign wireOut[185] = wireIn[186];    
  assign wireOut[186] = wireIn[185];    
  assign wireOut[187] = wireIn[187];    
  assign wireOut[188] = wireIn[188];    
  assign wireOut[189] = wireIn[190];    
  assign wireOut[190] = wireIn[189];    
  assign wireOut[191] = wireIn[191];    
  assign wireOut[192] = wireIn[192];    
  assign wireOut[193] = wireIn[194];    
  assign wireOut[194] = wireIn[193];    
  assign wireOut[195] = wireIn[195];    
  assign wireOut[196] = wireIn[196];    
  assign wireOut[197] = wireIn[198];    
  assign wireOut[198] = wireIn[197];    
  assign wireOut[199] = wireIn[199];    
  assign wireOut[200] = wireIn[200];    
  assign wireOut[201] = wireIn[202];    
  assign wireOut[202] = wireIn[201];    
  assign wireOut[203] = wireIn[203];    
  assign wireOut[204] = wireIn[204];    
  assign wireOut[205] = wireIn[206];    
  assign wireOut[206] = wireIn[205];    
  assign wireOut[207] = wireIn[207];    
  assign wireOut[208] = wireIn[208];    
  assign wireOut[209] = wireIn[210];    
  assign wireOut[210] = wireIn[209];    
  assign wireOut[211] = wireIn[211];    
  assign wireOut[212] = wireIn[212];    
  assign wireOut[213] = wireIn[214];    
  assign wireOut[214] = wireIn[213];    
  assign wireOut[215] = wireIn[215];    
  assign wireOut[216] = wireIn[216];    
  assign wireOut[217] = wireIn[218];    
  assign wireOut[218] = wireIn[217];    
  assign wireOut[219] = wireIn[219];    
  assign wireOut[220] = wireIn[220];    
  assign wireOut[221] = wireIn[222];    
  assign wireOut[222] = wireIn[221];    
  assign wireOut[223] = wireIn[223];    
  assign wireOut[224] = wireIn[224];    
  assign wireOut[225] = wireIn[226];    
  assign wireOut[226] = wireIn[225];    
  assign wireOut[227] = wireIn[227];    
  assign wireOut[228] = wireIn[228];    
  assign wireOut[229] = wireIn[230];    
  assign wireOut[230] = wireIn[229];    
  assign wireOut[231] = wireIn[231];    
  assign wireOut[232] = wireIn[232];    
  assign wireOut[233] = wireIn[234];    
  assign wireOut[234] = wireIn[233];    
  assign wireOut[235] = wireIn[235];    
  assign wireOut[236] = wireIn[236];    
  assign wireOut[237] = wireIn[238];    
  assign wireOut[238] = wireIn[237];    
  assign wireOut[239] = wireIn[239];    
  assign wireOut[240] = wireIn[240];    
  assign wireOut[241] = wireIn[242];    
  assign wireOut[242] = wireIn[241];    
  assign wireOut[243] = wireIn[243];    
  assign wireOut[244] = wireIn[244];    
  assign wireOut[245] = wireIn[246];    
  assign wireOut[246] = wireIn[245];    
  assign wireOut[247] = wireIn[247];    
  assign wireOut[248] = wireIn[248];    
  assign wireOut[249] = wireIn[250];    
  assign wireOut[250] = wireIn[249];    
  assign wireOut[251] = wireIn[251];    
  assign wireOut[252] = wireIn[252];    
  assign wireOut[253] = wireIn[254];    
  assign wireOut[254] = wireIn[253];    
  assign wireOut[255] = wireIn[255];    
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module switches_stage_st7_0_R(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
ctrl,                            
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;                   
  input [128-1:0] ctrl;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  switch_2_2 switch_inst_0(.inData_0(wireIn[0]), .inData_1(wireIn[1]), .outData_0(wireOut[0]), .outData_1(wireOut[1]), .ctrl(ctrl[0]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_1(.inData_0(wireIn[2]), .inData_1(wireIn[3]), .outData_0(wireOut[2]), .outData_1(wireOut[3]), .ctrl(ctrl[1]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_2(.inData_0(wireIn[4]), .inData_1(wireIn[5]), .outData_0(wireOut[4]), .outData_1(wireOut[5]), .ctrl(ctrl[2]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_3(.inData_0(wireIn[6]), .inData_1(wireIn[7]), .outData_0(wireOut[6]), .outData_1(wireOut[7]), .ctrl(ctrl[3]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_4(.inData_0(wireIn[8]), .inData_1(wireIn[9]), .outData_0(wireOut[8]), .outData_1(wireOut[9]), .ctrl(ctrl[4]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_5(.inData_0(wireIn[10]), .inData_1(wireIn[11]), .outData_0(wireOut[10]), .outData_1(wireOut[11]), .ctrl(ctrl[5]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_6(.inData_0(wireIn[12]), .inData_1(wireIn[13]), .outData_0(wireOut[12]), .outData_1(wireOut[13]), .ctrl(ctrl[6]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_7(.inData_0(wireIn[14]), .inData_1(wireIn[15]), .outData_0(wireOut[14]), .outData_1(wireOut[15]), .ctrl(ctrl[7]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_8(.inData_0(wireIn[16]), .inData_1(wireIn[17]), .outData_0(wireOut[16]), .outData_1(wireOut[17]), .ctrl(ctrl[8]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_9(.inData_0(wireIn[18]), .inData_1(wireIn[19]), .outData_0(wireOut[18]), .outData_1(wireOut[19]), .ctrl(ctrl[9]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_10(.inData_0(wireIn[20]), .inData_1(wireIn[21]), .outData_0(wireOut[20]), .outData_1(wireOut[21]), .ctrl(ctrl[10]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_11(.inData_0(wireIn[22]), .inData_1(wireIn[23]), .outData_0(wireOut[22]), .outData_1(wireOut[23]), .ctrl(ctrl[11]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_12(.inData_0(wireIn[24]), .inData_1(wireIn[25]), .outData_0(wireOut[24]), .outData_1(wireOut[25]), .ctrl(ctrl[12]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_13(.inData_0(wireIn[26]), .inData_1(wireIn[27]), .outData_0(wireOut[26]), .outData_1(wireOut[27]), .ctrl(ctrl[13]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_14(.inData_0(wireIn[28]), .inData_1(wireIn[29]), .outData_0(wireOut[28]), .outData_1(wireOut[29]), .ctrl(ctrl[14]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_15(.inData_0(wireIn[30]), .inData_1(wireIn[31]), .outData_0(wireOut[30]), .outData_1(wireOut[31]), .ctrl(ctrl[15]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_16(.inData_0(wireIn[32]), .inData_1(wireIn[33]), .outData_0(wireOut[32]), .outData_1(wireOut[33]), .ctrl(ctrl[16]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_17(.inData_0(wireIn[34]), .inData_1(wireIn[35]), .outData_0(wireOut[34]), .outData_1(wireOut[35]), .ctrl(ctrl[17]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_18(.inData_0(wireIn[36]), .inData_1(wireIn[37]), .outData_0(wireOut[36]), .outData_1(wireOut[37]), .ctrl(ctrl[18]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_19(.inData_0(wireIn[38]), .inData_1(wireIn[39]), .outData_0(wireOut[38]), .outData_1(wireOut[39]), .ctrl(ctrl[19]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_20(.inData_0(wireIn[40]), .inData_1(wireIn[41]), .outData_0(wireOut[40]), .outData_1(wireOut[41]), .ctrl(ctrl[20]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_21(.inData_0(wireIn[42]), .inData_1(wireIn[43]), .outData_0(wireOut[42]), .outData_1(wireOut[43]), .ctrl(ctrl[21]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_22(.inData_0(wireIn[44]), .inData_1(wireIn[45]), .outData_0(wireOut[44]), .outData_1(wireOut[45]), .ctrl(ctrl[22]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_23(.inData_0(wireIn[46]), .inData_1(wireIn[47]), .outData_0(wireOut[46]), .outData_1(wireOut[47]), .ctrl(ctrl[23]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_24(.inData_0(wireIn[48]), .inData_1(wireIn[49]), .outData_0(wireOut[48]), .outData_1(wireOut[49]), .ctrl(ctrl[24]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_25(.inData_0(wireIn[50]), .inData_1(wireIn[51]), .outData_0(wireOut[50]), .outData_1(wireOut[51]), .ctrl(ctrl[25]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_26(.inData_0(wireIn[52]), .inData_1(wireIn[53]), .outData_0(wireOut[52]), .outData_1(wireOut[53]), .ctrl(ctrl[26]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_27(.inData_0(wireIn[54]), .inData_1(wireIn[55]), .outData_0(wireOut[54]), .outData_1(wireOut[55]), .ctrl(ctrl[27]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_28(.inData_0(wireIn[56]), .inData_1(wireIn[57]), .outData_0(wireOut[56]), .outData_1(wireOut[57]), .ctrl(ctrl[28]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_29(.inData_0(wireIn[58]), .inData_1(wireIn[59]), .outData_0(wireOut[58]), .outData_1(wireOut[59]), .ctrl(ctrl[29]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_30(.inData_0(wireIn[60]), .inData_1(wireIn[61]), .outData_0(wireOut[60]), .outData_1(wireOut[61]), .ctrl(ctrl[30]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_31(.inData_0(wireIn[62]), .inData_1(wireIn[63]), .outData_0(wireOut[62]), .outData_1(wireOut[63]), .ctrl(ctrl[31]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_32(.inData_0(wireIn[64]), .inData_1(wireIn[65]), .outData_0(wireOut[64]), .outData_1(wireOut[65]), .ctrl(ctrl[32]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_33(.inData_0(wireIn[66]), .inData_1(wireIn[67]), .outData_0(wireOut[66]), .outData_1(wireOut[67]), .ctrl(ctrl[33]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_34(.inData_0(wireIn[68]), .inData_1(wireIn[69]), .outData_0(wireOut[68]), .outData_1(wireOut[69]), .ctrl(ctrl[34]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_35(.inData_0(wireIn[70]), .inData_1(wireIn[71]), .outData_0(wireOut[70]), .outData_1(wireOut[71]), .ctrl(ctrl[35]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_36(.inData_0(wireIn[72]), .inData_1(wireIn[73]), .outData_0(wireOut[72]), .outData_1(wireOut[73]), .ctrl(ctrl[36]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_37(.inData_0(wireIn[74]), .inData_1(wireIn[75]), .outData_0(wireOut[74]), .outData_1(wireOut[75]), .ctrl(ctrl[37]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_38(.inData_0(wireIn[76]), .inData_1(wireIn[77]), .outData_0(wireOut[76]), .outData_1(wireOut[77]), .ctrl(ctrl[38]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_39(.inData_0(wireIn[78]), .inData_1(wireIn[79]), .outData_0(wireOut[78]), .outData_1(wireOut[79]), .ctrl(ctrl[39]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_40(.inData_0(wireIn[80]), .inData_1(wireIn[81]), .outData_0(wireOut[80]), .outData_1(wireOut[81]), .ctrl(ctrl[40]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_41(.inData_0(wireIn[82]), .inData_1(wireIn[83]), .outData_0(wireOut[82]), .outData_1(wireOut[83]), .ctrl(ctrl[41]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_42(.inData_0(wireIn[84]), .inData_1(wireIn[85]), .outData_0(wireOut[84]), .outData_1(wireOut[85]), .ctrl(ctrl[42]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_43(.inData_0(wireIn[86]), .inData_1(wireIn[87]), .outData_0(wireOut[86]), .outData_1(wireOut[87]), .ctrl(ctrl[43]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_44(.inData_0(wireIn[88]), .inData_1(wireIn[89]), .outData_0(wireOut[88]), .outData_1(wireOut[89]), .ctrl(ctrl[44]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_45(.inData_0(wireIn[90]), .inData_1(wireIn[91]), .outData_0(wireOut[90]), .outData_1(wireOut[91]), .ctrl(ctrl[45]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_46(.inData_0(wireIn[92]), .inData_1(wireIn[93]), .outData_0(wireOut[92]), .outData_1(wireOut[93]), .ctrl(ctrl[46]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_47(.inData_0(wireIn[94]), .inData_1(wireIn[95]), .outData_0(wireOut[94]), .outData_1(wireOut[95]), .ctrl(ctrl[47]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_48(.inData_0(wireIn[96]), .inData_1(wireIn[97]), .outData_0(wireOut[96]), .outData_1(wireOut[97]), .ctrl(ctrl[48]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_49(.inData_0(wireIn[98]), .inData_1(wireIn[99]), .outData_0(wireOut[98]), .outData_1(wireOut[99]), .ctrl(ctrl[49]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_50(.inData_0(wireIn[100]), .inData_1(wireIn[101]), .outData_0(wireOut[100]), .outData_1(wireOut[101]), .ctrl(ctrl[50]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_51(.inData_0(wireIn[102]), .inData_1(wireIn[103]), .outData_0(wireOut[102]), .outData_1(wireOut[103]), .ctrl(ctrl[51]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_52(.inData_0(wireIn[104]), .inData_1(wireIn[105]), .outData_0(wireOut[104]), .outData_1(wireOut[105]), .ctrl(ctrl[52]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_53(.inData_0(wireIn[106]), .inData_1(wireIn[107]), .outData_0(wireOut[106]), .outData_1(wireOut[107]), .ctrl(ctrl[53]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_54(.inData_0(wireIn[108]), .inData_1(wireIn[109]), .outData_0(wireOut[108]), .outData_1(wireOut[109]), .ctrl(ctrl[54]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_55(.inData_0(wireIn[110]), .inData_1(wireIn[111]), .outData_0(wireOut[110]), .outData_1(wireOut[111]), .ctrl(ctrl[55]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_56(.inData_0(wireIn[112]), .inData_1(wireIn[113]), .outData_0(wireOut[112]), .outData_1(wireOut[113]), .ctrl(ctrl[56]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_57(.inData_0(wireIn[114]), .inData_1(wireIn[115]), .outData_0(wireOut[114]), .outData_1(wireOut[115]), .ctrl(ctrl[57]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_58(.inData_0(wireIn[116]), .inData_1(wireIn[117]), .outData_0(wireOut[116]), .outData_1(wireOut[117]), .ctrl(ctrl[58]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_59(.inData_0(wireIn[118]), .inData_1(wireIn[119]), .outData_0(wireOut[118]), .outData_1(wireOut[119]), .ctrl(ctrl[59]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_60(.inData_0(wireIn[120]), .inData_1(wireIn[121]), .outData_0(wireOut[120]), .outData_1(wireOut[121]), .ctrl(ctrl[60]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_61(.inData_0(wireIn[122]), .inData_1(wireIn[123]), .outData_0(wireOut[122]), .outData_1(wireOut[123]), .ctrl(ctrl[61]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_62(.inData_0(wireIn[124]), .inData_1(wireIn[125]), .outData_0(wireOut[124]), .outData_1(wireOut[125]), .ctrl(ctrl[62]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_63(.inData_0(wireIn[126]), .inData_1(wireIn[127]), .outData_0(wireOut[126]), .outData_1(wireOut[127]), .ctrl(ctrl[63]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_64(.inData_0(wireIn[128]), .inData_1(wireIn[129]), .outData_0(wireOut[128]), .outData_1(wireOut[129]), .ctrl(ctrl[64]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_65(.inData_0(wireIn[130]), .inData_1(wireIn[131]), .outData_0(wireOut[130]), .outData_1(wireOut[131]), .ctrl(ctrl[65]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_66(.inData_0(wireIn[132]), .inData_1(wireIn[133]), .outData_0(wireOut[132]), .outData_1(wireOut[133]), .ctrl(ctrl[66]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_67(.inData_0(wireIn[134]), .inData_1(wireIn[135]), .outData_0(wireOut[134]), .outData_1(wireOut[135]), .ctrl(ctrl[67]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_68(.inData_0(wireIn[136]), .inData_1(wireIn[137]), .outData_0(wireOut[136]), .outData_1(wireOut[137]), .ctrl(ctrl[68]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_69(.inData_0(wireIn[138]), .inData_1(wireIn[139]), .outData_0(wireOut[138]), .outData_1(wireOut[139]), .ctrl(ctrl[69]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_70(.inData_0(wireIn[140]), .inData_1(wireIn[141]), .outData_0(wireOut[140]), .outData_1(wireOut[141]), .ctrl(ctrl[70]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_71(.inData_0(wireIn[142]), .inData_1(wireIn[143]), .outData_0(wireOut[142]), .outData_1(wireOut[143]), .ctrl(ctrl[71]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_72(.inData_0(wireIn[144]), .inData_1(wireIn[145]), .outData_0(wireOut[144]), .outData_1(wireOut[145]), .ctrl(ctrl[72]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_73(.inData_0(wireIn[146]), .inData_1(wireIn[147]), .outData_0(wireOut[146]), .outData_1(wireOut[147]), .ctrl(ctrl[73]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_74(.inData_0(wireIn[148]), .inData_1(wireIn[149]), .outData_0(wireOut[148]), .outData_1(wireOut[149]), .ctrl(ctrl[74]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_75(.inData_0(wireIn[150]), .inData_1(wireIn[151]), .outData_0(wireOut[150]), .outData_1(wireOut[151]), .ctrl(ctrl[75]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_76(.inData_0(wireIn[152]), .inData_1(wireIn[153]), .outData_0(wireOut[152]), .outData_1(wireOut[153]), .ctrl(ctrl[76]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_77(.inData_0(wireIn[154]), .inData_1(wireIn[155]), .outData_0(wireOut[154]), .outData_1(wireOut[155]), .ctrl(ctrl[77]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_78(.inData_0(wireIn[156]), .inData_1(wireIn[157]), .outData_0(wireOut[156]), .outData_1(wireOut[157]), .ctrl(ctrl[78]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_79(.inData_0(wireIn[158]), .inData_1(wireIn[159]), .outData_0(wireOut[158]), .outData_1(wireOut[159]), .ctrl(ctrl[79]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_80(.inData_0(wireIn[160]), .inData_1(wireIn[161]), .outData_0(wireOut[160]), .outData_1(wireOut[161]), .ctrl(ctrl[80]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_81(.inData_0(wireIn[162]), .inData_1(wireIn[163]), .outData_0(wireOut[162]), .outData_1(wireOut[163]), .ctrl(ctrl[81]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_82(.inData_0(wireIn[164]), .inData_1(wireIn[165]), .outData_0(wireOut[164]), .outData_1(wireOut[165]), .ctrl(ctrl[82]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_83(.inData_0(wireIn[166]), .inData_1(wireIn[167]), .outData_0(wireOut[166]), .outData_1(wireOut[167]), .ctrl(ctrl[83]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_84(.inData_0(wireIn[168]), .inData_1(wireIn[169]), .outData_0(wireOut[168]), .outData_1(wireOut[169]), .ctrl(ctrl[84]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_85(.inData_0(wireIn[170]), .inData_1(wireIn[171]), .outData_0(wireOut[170]), .outData_1(wireOut[171]), .ctrl(ctrl[85]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_86(.inData_0(wireIn[172]), .inData_1(wireIn[173]), .outData_0(wireOut[172]), .outData_1(wireOut[173]), .ctrl(ctrl[86]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_87(.inData_0(wireIn[174]), .inData_1(wireIn[175]), .outData_0(wireOut[174]), .outData_1(wireOut[175]), .ctrl(ctrl[87]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_88(.inData_0(wireIn[176]), .inData_1(wireIn[177]), .outData_0(wireOut[176]), .outData_1(wireOut[177]), .ctrl(ctrl[88]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_89(.inData_0(wireIn[178]), .inData_1(wireIn[179]), .outData_0(wireOut[178]), .outData_1(wireOut[179]), .ctrl(ctrl[89]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_90(.inData_0(wireIn[180]), .inData_1(wireIn[181]), .outData_0(wireOut[180]), .outData_1(wireOut[181]), .ctrl(ctrl[90]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_91(.inData_0(wireIn[182]), .inData_1(wireIn[183]), .outData_0(wireOut[182]), .outData_1(wireOut[183]), .ctrl(ctrl[91]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_92(.inData_0(wireIn[184]), .inData_1(wireIn[185]), .outData_0(wireOut[184]), .outData_1(wireOut[185]), .ctrl(ctrl[92]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_93(.inData_0(wireIn[186]), .inData_1(wireIn[187]), .outData_0(wireOut[186]), .outData_1(wireOut[187]), .ctrl(ctrl[93]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_94(.inData_0(wireIn[188]), .inData_1(wireIn[189]), .outData_0(wireOut[188]), .outData_1(wireOut[189]), .ctrl(ctrl[94]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_95(.inData_0(wireIn[190]), .inData_1(wireIn[191]), .outData_0(wireOut[190]), .outData_1(wireOut[191]), .ctrl(ctrl[95]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_96(.inData_0(wireIn[192]), .inData_1(wireIn[193]), .outData_0(wireOut[192]), .outData_1(wireOut[193]), .ctrl(ctrl[96]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_97(.inData_0(wireIn[194]), .inData_1(wireIn[195]), .outData_0(wireOut[194]), .outData_1(wireOut[195]), .ctrl(ctrl[97]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_98(.inData_0(wireIn[196]), .inData_1(wireIn[197]), .outData_0(wireOut[196]), .outData_1(wireOut[197]), .ctrl(ctrl[98]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_99(.inData_0(wireIn[198]), .inData_1(wireIn[199]), .outData_0(wireOut[198]), .outData_1(wireOut[199]), .ctrl(ctrl[99]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_100(.inData_0(wireIn[200]), .inData_1(wireIn[201]), .outData_0(wireOut[200]), .outData_1(wireOut[201]), .ctrl(ctrl[100]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_101(.inData_0(wireIn[202]), .inData_1(wireIn[203]), .outData_0(wireOut[202]), .outData_1(wireOut[203]), .ctrl(ctrl[101]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_102(.inData_0(wireIn[204]), .inData_1(wireIn[205]), .outData_0(wireOut[204]), .outData_1(wireOut[205]), .ctrl(ctrl[102]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_103(.inData_0(wireIn[206]), .inData_1(wireIn[207]), .outData_0(wireOut[206]), .outData_1(wireOut[207]), .ctrl(ctrl[103]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_104(.inData_0(wireIn[208]), .inData_1(wireIn[209]), .outData_0(wireOut[208]), .outData_1(wireOut[209]), .ctrl(ctrl[104]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_105(.inData_0(wireIn[210]), .inData_1(wireIn[211]), .outData_0(wireOut[210]), .outData_1(wireOut[211]), .ctrl(ctrl[105]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_106(.inData_0(wireIn[212]), .inData_1(wireIn[213]), .outData_0(wireOut[212]), .outData_1(wireOut[213]), .ctrl(ctrl[106]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_107(.inData_0(wireIn[214]), .inData_1(wireIn[215]), .outData_0(wireOut[214]), .outData_1(wireOut[215]), .ctrl(ctrl[107]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_108(.inData_0(wireIn[216]), .inData_1(wireIn[217]), .outData_0(wireOut[216]), .outData_1(wireOut[217]), .ctrl(ctrl[108]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_109(.inData_0(wireIn[218]), .inData_1(wireIn[219]), .outData_0(wireOut[218]), .outData_1(wireOut[219]), .ctrl(ctrl[109]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_110(.inData_0(wireIn[220]), .inData_1(wireIn[221]), .outData_0(wireOut[220]), .outData_1(wireOut[221]), .ctrl(ctrl[110]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_111(.inData_0(wireIn[222]), .inData_1(wireIn[223]), .outData_0(wireOut[222]), .outData_1(wireOut[223]), .ctrl(ctrl[111]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_112(.inData_0(wireIn[224]), .inData_1(wireIn[225]), .outData_0(wireOut[224]), .outData_1(wireOut[225]), .ctrl(ctrl[112]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_113(.inData_0(wireIn[226]), .inData_1(wireIn[227]), .outData_0(wireOut[226]), .outData_1(wireOut[227]), .ctrl(ctrl[113]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_114(.inData_0(wireIn[228]), .inData_1(wireIn[229]), .outData_0(wireOut[228]), .outData_1(wireOut[229]), .ctrl(ctrl[114]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_115(.inData_0(wireIn[230]), .inData_1(wireIn[231]), .outData_0(wireOut[230]), .outData_1(wireOut[231]), .ctrl(ctrl[115]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_116(.inData_0(wireIn[232]), .inData_1(wireIn[233]), .outData_0(wireOut[232]), .outData_1(wireOut[233]), .ctrl(ctrl[116]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_117(.inData_0(wireIn[234]), .inData_1(wireIn[235]), .outData_0(wireOut[234]), .outData_1(wireOut[235]), .ctrl(ctrl[117]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_118(.inData_0(wireIn[236]), .inData_1(wireIn[237]), .outData_0(wireOut[236]), .outData_1(wireOut[237]), .ctrl(ctrl[118]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_119(.inData_0(wireIn[238]), .inData_1(wireIn[239]), .outData_0(wireOut[238]), .outData_1(wireOut[239]), .ctrl(ctrl[119]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_120(.inData_0(wireIn[240]), .inData_1(wireIn[241]), .outData_0(wireOut[240]), .outData_1(wireOut[241]), .ctrl(ctrl[120]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_121(.inData_0(wireIn[242]), .inData_1(wireIn[243]), .outData_0(wireOut[242]), .outData_1(wireOut[243]), .ctrl(ctrl[121]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_122(.inData_0(wireIn[244]), .inData_1(wireIn[245]), .outData_0(wireOut[244]), .outData_1(wireOut[245]), .ctrl(ctrl[122]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_123(.inData_0(wireIn[246]), .inData_1(wireIn[247]), .outData_0(wireOut[246]), .outData_1(wireOut[247]), .ctrl(ctrl[123]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_124(.inData_0(wireIn[248]), .inData_1(wireIn[249]), .outData_0(wireOut[248]), .outData_1(wireOut[249]), .ctrl(ctrl[124]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_125(.inData_0(wireIn[250]), .inData_1(wireIn[251]), .outData_0(wireOut[250]), .outData_1(wireOut[251]), .ctrl(ctrl[125]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_126(.inData_0(wireIn[252]), .inData_1(wireIn[253]), .outData_0(wireOut[252]), .outData_1(wireOut[253]), .ctrl(ctrl[126]), .clk(clk), .rst(rst));
  switch_2_2 switch_inst_127(.inData_0(wireIn[254]), .inData_1(wireIn[255]), .outData_0(wireOut[254]), .outData_1(wireOut[255]), .ctrl(ctrl[127]), .clk(clk), .rst(rst));
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module wireCon_dp256_st7_R(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  assign wireOut[0] = wireIn[0];    
  assign wireOut[1] = wireIn[1];    
  assign wireOut[2] = wireIn[2];    
  assign wireOut[3] = wireIn[3];    
  assign wireOut[4] = wireIn[4];    
  assign wireOut[5] = wireIn[5];    
  assign wireOut[6] = wireIn[6];    
  assign wireOut[7] = wireIn[7];    
  assign wireOut[8] = wireIn[8];    
  assign wireOut[9] = wireIn[9];    
  assign wireOut[10] = wireIn[10];    
  assign wireOut[11] = wireIn[11];    
  assign wireOut[12] = wireIn[12];    
  assign wireOut[13] = wireIn[13];    
  assign wireOut[14] = wireIn[14];    
  assign wireOut[15] = wireIn[15];    
  assign wireOut[16] = wireIn[16];    
  assign wireOut[17] = wireIn[17];    
  assign wireOut[18] = wireIn[18];    
  assign wireOut[19] = wireIn[19];    
  assign wireOut[20] = wireIn[20];    
  assign wireOut[21] = wireIn[21];    
  assign wireOut[22] = wireIn[22];    
  assign wireOut[23] = wireIn[23];    
  assign wireOut[24] = wireIn[24];    
  assign wireOut[25] = wireIn[25];    
  assign wireOut[26] = wireIn[26];    
  assign wireOut[27] = wireIn[27];    
  assign wireOut[28] = wireIn[28];    
  assign wireOut[29] = wireIn[29];    
  assign wireOut[30] = wireIn[30];    
  assign wireOut[31] = wireIn[31];    
  assign wireOut[32] = wireIn[32];    
  assign wireOut[33] = wireIn[33];    
  assign wireOut[34] = wireIn[34];    
  assign wireOut[35] = wireIn[35];    
  assign wireOut[36] = wireIn[36];    
  assign wireOut[37] = wireIn[37];    
  assign wireOut[38] = wireIn[38];    
  assign wireOut[39] = wireIn[39];    
  assign wireOut[40] = wireIn[40];    
  assign wireOut[41] = wireIn[41];    
  assign wireOut[42] = wireIn[42];    
  assign wireOut[43] = wireIn[43];    
  assign wireOut[44] = wireIn[44];    
  assign wireOut[45] = wireIn[45];    
  assign wireOut[46] = wireIn[46];    
  assign wireOut[47] = wireIn[47];    
  assign wireOut[48] = wireIn[48];    
  assign wireOut[49] = wireIn[49];    
  assign wireOut[50] = wireIn[50];    
  assign wireOut[51] = wireIn[51];    
  assign wireOut[52] = wireIn[52];    
  assign wireOut[53] = wireIn[53];    
  assign wireOut[54] = wireIn[54];    
  assign wireOut[55] = wireIn[55];    
  assign wireOut[56] = wireIn[56];    
  assign wireOut[57] = wireIn[57];    
  assign wireOut[58] = wireIn[58];    
  assign wireOut[59] = wireIn[59];    
  assign wireOut[60] = wireIn[60];    
  assign wireOut[61] = wireIn[61];    
  assign wireOut[62] = wireIn[62];    
  assign wireOut[63] = wireIn[63];    
  assign wireOut[64] = wireIn[64];    
  assign wireOut[65] = wireIn[65];    
  assign wireOut[66] = wireIn[66];    
  assign wireOut[67] = wireIn[67];    
  assign wireOut[68] = wireIn[68];    
  assign wireOut[69] = wireIn[69];    
  assign wireOut[70] = wireIn[70];    
  assign wireOut[71] = wireIn[71];    
  assign wireOut[72] = wireIn[72];    
  assign wireOut[73] = wireIn[73];    
  assign wireOut[74] = wireIn[74];    
  assign wireOut[75] = wireIn[75];    
  assign wireOut[76] = wireIn[76];    
  assign wireOut[77] = wireIn[77];    
  assign wireOut[78] = wireIn[78];    
  assign wireOut[79] = wireIn[79];    
  assign wireOut[80] = wireIn[80];    
  assign wireOut[81] = wireIn[81];    
  assign wireOut[82] = wireIn[82];    
  assign wireOut[83] = wireIn[83];    
  assign wireOut[84] = wireIn[84];    
  assign wireOut[85] = wireIn[85];    
  assign wireOut[86] = wireIn[86];    
  assign wireOut[87] = wireIn[87];    
  assign wireOut[88] = wireIn[88];    
  assign wireOut[89] = wireIn[89];    
  assign wireOut[90] = wireIn[90];    
  assign wireOut[91] = wireIn[91];    
  assign wireOut[92] = wireIn[92];    
  assign wireOut[93] = wireIn[93];    
  assign wireOut[94] = wireIn[94];    
  assign wireOut[95] = wireIn[95];    
  assign wireOut[96] = wireIn[96];    
  assign wireOut[97] = wireIn[97];    
  assign wireOut[98] = wireIn[98];    
  assign wireOut[99] = wireIn[99];    
  assign wireOut[100] = wireIn[100];    
  assign wireOut[101] = wireIn[101];    
  assign wireOut[102] = wireIn[102];    
  assign wireOut[103] = wireIn[103];    
  assign wireOut[104] = wireIn[104];    
  assign wireOut[105] = wireIn[105];    
  assign wireOut[106] = wireIn[106];    
  assign wireOut[107] = wireIn[107];    
  assign wireOut[108] = wireIn[108];    
  assign wireOut[109] = wireIn[109];    
  assign wireOut[110] = wireIn[110];    
  assign wireOut[111] = wireIn[111];    
  assign wireOut[112] = wireIn[112];    
  assign wireOut[113] = wireIn[113];    
  assign wireOut[114] = wireIn[114];    
  assign wireOut[115] = wireIn[115];    
  assign wireOut[116] = wireIn[116];    
  assign wireOut[117] = wireIn[117];    
  assign wireOut[118] = wireIn[118];    
  assign wireOut[119] = wireIn[119];    
  assign wireOut[120] = wireIn[120];    
  assign wireOut[121] = wireIn[121];    
  assign wireOut[122] = wireIn[122];    
  assign wireOut[123] = wireIn[123];    
  assign wireOut[124] = wireIn[124];    
  assign wireOut[125] = wireIn[125];    
  assign wireOut[126] = wireIn[126];    
  assign wireOut[127] = wireIn[127];    
  assign wireOut[128] = wireIn[128];    
  assign wireOut[129] = wireIn[129];    
  assign wireOut[130] = wireIn[130];    
  assign wireOut[131] = wireIn[131];    
  assign wireOut[132] = wireIn[132];    
  assign wireOut[133] = wireIn[133];    
  assign wireOut[134] = wireIn[134];    
  assign wireOut[135] = wireIn[135];    
  assign wireOut[136] = wireIn[136];    
  assign wireOut[137] = wireIn[137];    
  assign wireOut[138] = wireIn[138];    
  assign wireOut[139] = wireIn[139];    
  assign wireOut[140] = wireIn[140];    
  assign wireOut[141] = wireIn[141];    
  assign wireOut[142] = wireIn[142];    
  assign wireOut[143] = wireIn[143];    
  assign wireOut[144] = wireIn[144];    
  assign wireOut[145] = wireIn[145];    
  assign wireOut[146] = wireIn[146];    
  assign wireOut[147] = wireIn[147];    
  assign wireOut[148] = wireIn[148];    
  assign wireOut[149] = wireIn[149];    
  assign wireOut[150] = wireIn[150];    
  assign wireOut[151] = wireIn[151];    
  assign wireOut[152] = wireIn[152];    
  assign wireOut[153] = wireIn[153];    
  assign wireOut[154] = wireIn[154];    
  assign wireOut[155] = wireIn[155];    
  assign wireOut[156] = wireIn[156];    
  assign wireOut[157] = wireIn[157];    
  assign wireOut[158] = wireIn[158];    
  assign wireOut[159] = wireIn[159];    
  assign wireOut[160] = wireIn[160];    
  assign wireOut[161] = wireIn[161];    
  assign wireOut[162] = wireIn[162];    
  assign wireOut[163] = wireIn[163];    
  assign wireOut[164] = wireIn[164];    
  assign wireOut[165] = wireIn[165];    
  assign wireOut[166] = wireIn[166];    
  assign wireOut[167] = wireIn[167];    
  assign wireOut[168] = wireIn[168];    
  assign wireOut[169] = wireIn[169];    
  assign wireOut[170] = wireIn[170];    
  assign wireOut[171] = wireIn[171];    
  assign wireOut[172] = wireIn[172];    
  assign wireOut[173] = wireIn[173];    
  assign wireOut[174] = wireIn[174];    
  assign wireOut[175] = wireIn[175];    
  assign wireOut[176] = wireIn[176];    
  assign wireOut[177] = wireIn[177];    
  assign wireOut[178] = wireIn[178];    
  assign wireOut[179] = wireIn[179];    
  assign wireOut[180] = wireIn[180];    
  assign wireOut[181] = wireIn[181];    
  assign wireOut[182] = wireIn[182];    
  assign wireOut[183] = wireIn[183];    
  assign wireOut[184] = wireIn[184];    
  assign wireOut[185] = wireIn[185];    
  assign wireOut[186] = wireIn[186];    
  assign wireOut[187] = wireIn[187];    
  assign wireOut[188] = wireIn[188];    
  assign wireOut[189] = wireIn[189];    
  assign wireOut[190] = wireIn[190];    
  assign wireOut[191] = wireIn[191];    
  assign wireOut[192] = wireIn[192];    
  assign wireOut[193] = wireIn[193];    
  assign wireOut[194] = wireIn[194];    
  assign wireOut[195] = wireIn[195];    
  assign wireOut[196] = wireIn[196];    
  assign wireOut[197] = wireIn[197];    
  assign wireOut[198] = wireIn[198];    
  assign wireOut[199] = wireIn[199];    
  assign wireOut[200] = wireIn[200];    
  assign wireOut[201] = wireIn[201];    
  assign wireOut[202] = wireIn[202];    
  assign wireOut[203] = wireIn[203];    
  assign wireOut[204] = wireIn[204];    
  assign wireOut[205] = wireIn[205];    
  assign wireOut[206] = wireIn[206];    
  assign wireOut[207] = wireIn[207];    
  assign wireOut[208] = wireIn[208];    
  assign wireOut[209] = wireIn[209];    
  assign wireOut[210] = wireIn[210];    
  assign wireOut[211] = wireIn[211];    
  assign wireOut[212] = wireIn[212];    
  assign wireOut[213] = wireIn[213];    
  assign wireOut[214] = wireIn[214];    
  assign wireOut[215] = wireIn[215];    
  assign wireOut[216] = wireIn[216];    
  assign wireOut[217] = wireIn[217];    
  assign wireOut[218] = wireIn[218];    
  assign wireOut[219] = wireIn[219];    
  assign wireOut[220] = wireIn[220];    
  assign wireOut[221] = wireIn[221];    
  assign wireOut[222] = wireIn[222];    
  assign wireOut[223] = wireIn[223];    
  assign wireOut[224] = wireIn[224];    
  assign wireOut[225] = wireIn[225];    
  assign wireOut[226] = wireIn[226];    
  assign wireOut[227] = wireIn[227];    
  assign wireOut[228] = wireIn[228];    
  assign wireOut[229] = wireIn[229];    
  assign wireOut[230] = wireIn[230];    
  assign wireOut[231] = wireIn[231];    
  assign wireOut[232] = wireIn[232];    
  assign wireOut[233] = wireIn[233];    
  assign wireOut[234] = wireIn[234];    
  assign wireOut[235] = wireIn[235];    
  assign wireOut[236] = wireIn[236];    
  assign wireOut[237] = wireIn[237];    
  assign wireOut[238] = wireIn[238];    
  assign wireOut[239] = wireIn[239];    
  assign wireOut[240] = wireIn[240];    
  assign wireOut[241] = wireIn[241];    
  assign wireOut[242] = wireIn[242];    
  assign wireOut[243] = wireIn[243];    
  assign wireOut[244] = wireIn[244];    
  assign wireOut[245] = wireIn[245];    
  assign wireOut[246] = wireIn[246];    
  assign wireOut[247] = wireIn[247];    
  assign wireOut[248] = wireIn[248];    
  assign wireOut[249] = wireIn[249];    
  assign wireOut[250] = wireIn[250];    
  assign wireOut[251] = wireIn[251];    
  assign wireOut[252] = wireIn[252];    
  assign wireOut[253] = wireIn[253];    
  assign wireOut[254] = wireIn[254];    
  assign wireOut[255] = wireIn[255];    
  
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = in_start;    
  
endmodule                        


module egressStage_p256(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
counter_in,                       
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;                   
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  input [7:0] counter_in; 
  output [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255;
  output out_start; 
  
  
  wire out_start_w; 
  wire [DATA_WIDTH-1:0] wireIn [255:0];              
  wire [DATA_WIDTH-1:0] wireOut [255:0];              
  
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  wire in_start_stage7;
  wire con_in_start_stage7;

  wire in_start_stage6;
  wire con_in_start_stage6;

  wire in_start_stage5;
  wire con_in_start_stage5;

  wire in_start_stage4;
  wire con_in_start_stage4;

  wire in_start_stage3;
  wire con_in_start_stage3;

  wire in_start_stage2;
  wire con_in_start_stage2;

  wire in_start_stage1;
  wire con_in_start_stage1;

  wire in_start_stage0;
  wire con_in_start_stage0;

  wire [DATA_WIDTH-1:0] wire_switch_in_stage7[255:0];
  wire [DATA_WIDTH-1:0] wire_switch_out_stage7[255:0];
  reg [127:0] wire_ctrl_stage7;

  switches_stage_st7_0_R switch_stage_7(
        .inData_0(wire_switch_in_stage7[0]), .inData_1(wire_switch_in_stage7[1]), .inData_2(wire_switch_in_stage7[2]), .inData_3(wire_switch_in_stage7[3]), .inData_4(wire_switch_in_stage7[4]), .inData_5(wire_switch_in_stage7[5]), .inData_6(wire_switch_in_stage7[6]), .inData_7(wire_switch_in_stage7[7]), .inData_8(wire_switch_in_stage7[8]), .inData_9(wire_switch_in_stage7[9]), .inData_10(wire_switch_in_stage7[10]), .inData_11(wire_switch_in_stage7[11]), .inData_12(wire_switch_in_stage7[12]), .inData_13(wire_switch_in_stage7[13]), .inData_14(wire_switch_in_stage7[14]), .inData_15(wire_switch_in_stage7[15]), .inData_16(wire_switch_in_stage7[16]), .inData_17(wire_switch_in_stage7[17]), .inData_18(wire_switch_in_stage7[18]), .inData_19(wire_switch_in_stage7[19]), .inData_20(wire_switch_in_stage7[20]), .inData_21(wire_switch_in_stage7[21]), .inData_22(wire_switch_in_stage7[22]), .inData_23(wire_switch_in_stage7[23]), .inData_24(wire_switch_in_stage7[24]), .inData_25(wire_switch_in_stage7[25]), .inData_26(wire_switch_in_stage7[26]), .inData_27(wire_switch_in_stage7[27]), .inData_28(wire_switch_in_stage7[28]), .inData_29(wire_switch_in_stage7[29]), .inData_30(wire_switch_in_stage7[30]), .inData_31(wire_switch_in_stage7[31]), .inData_32(wire_switch_in_stage7[32]), .inData_33(wire_switch_in_stage7[33]), .inData_34(wire_switch_in_stage7[34]), .inData_35(wire_switch_in_stage7[35]), .inData_36(wire_switch_in_stage7[36]), .inData_37(wire_switch_in_stage7[37]), .inData_38(wire_switch_in_stage7[38]), .inData_39(wire_switch_in_stage7[39]), .inData_40(wire_switch_in_stage7[40]), .inData_41(wire_switch_in_stage7[41]), .inData_42(wire_switch_in_stage7[42]), .inData_43(wire_switch_in_stage7[43]), .inData_44(wire_switch_in_stage7[44]), .inData_45(wire_switch_in_stage7[45]), .inData_46(wire_switch_in_stage7[46]), .inData_47(wire_switch_in_stage7[47]), .inData_48(wire_switch_in_stage7[48]), .inData_49(wire_switch_in_stage7[49]), .inData_50(wire_switch_in_stage7[50]), .inData_51(wire_switch_in_stage7[51]), .inData_52(wire_switch_in_stage7[52]), .inData_53(wire_switch_in_stage7[53]), .inData_54(wire_switch_in_stage7[54]), .inData_55(wire_switch_in_stage7[55]), .inData_56(wire_switch_in_stage7[56]), .inData_57(wire_switch_in_stage7[57]), .inData_58(wire_switch_in_stage7[58]), .inData_59(wire_switch_in_stage7[59]), .inData_60(wire_switch_in_stage7[60]), .inData_61(wire_switch_in_stage7[61]), .inData_62(wire_switch_in_stage7[62]), .inData_63(wire_switch_in_stage7[63]), .inData_64(wire_switch_in_stage7[64]), .inData_65(wire_switch_in_stage7[65]), .inData_66(wire_switch_in_stage7[66]), .inData_67(wire_switch_in_stage7[67]), .inData_68(wire_switch_in_stage7[68]), .inData_69(wire_switch_in_stage7[69]), .inData_70(wire_switch_in_stage7[70]), .inData_71(wire_switch_in_stage7[71]), .inData_72(wire_switch_in_stage7[72]), .inData_73(wire_switch_in_stage7[73]), .inData_74(wire_switch_in_stage7[74]), .inData_75(wire_switch_in_stage7[75]), .inData_76(wire_switch_in_stage7[76]), .inData_77(wire_switch_in_stage7[77]), .inData_78(wire_switch_in_stage7[78]), .inData_79(wire_switch_in_stage7[79]), .inData_80(wire_switch_in_stage7[80]), .inData_81(wire_switch_in_stage7[81]), .inData_82(wire_switch_in_stage7[82]), .inData_83(wire_switch_in_stage7[83]), .inData_84(wire_switch_in_stage7[84]), .inData_85(wire_switch_in_stage7[85]), .inData_86(wire_switch_in_stage7[86]), .inData_87(wire_switch_in_stage7[87]), .inData_88(wire_switch_in_stage7[88]), .inData_89(wire_switch_in_stage7[89]), .inData_90(wire_switch_in_stage7[90]), .inData_91(wire_switch_in_stage7[91]), .inData_92(wire_switch_in_stage7[92]), .inData_93(wire_switch_in_stage7[93]), .inData_94(wire_switch_in_stage7[94]), .inData_95(wire_switch_in_stage7[95]), .inData_96(wire_switch_in_stage7[96]), .inData_97(wire_switch_in_stage7[97]), .inData_98(wire_switch_in_stage7[98]), .inData_99(wire_switch_in_stage7[99]), .inData_100(wire_switch_in_stage7[100]), .inData_101(wire_switch_in_stage7[101]), .inData_102(wire_switch_in_stage7[102]), .inData_103(wire_switch_in_stage7[103]), .inData_104(wire_switch_in_stage7[104]), .inData_105(wire_switch_in_stage7[105]), .inData_106(wire_switch_in_stage7[106]), .inData_107(wire_switch_in_stage7[107]), .inData_108(wire_switch_in_stage7[108]), .inData_109(wire_switch_in_stage7[109]), .inData_110(wire_switch_in_stage7[110]), .inData_111(wire_switch_in_stage7[111]), .inData_112(wire_switch_in_stage7[112]), .inData_113(wire_switch_in_stage7[113]), .inData_114(wire_switch_in_stage7[114]), .inData_115(wire_switch_in_stage7[115]), .inData_116(wire_switch_in_stage7[116]), .inData_117(wire_switch_in_stage7[117]), .inData_118(wire_switch_in_stage7[118]), .inData_119(wire_switch_in_stage7[119]), .inData_120(wire_switch_in_stage7[120]), .inData_121(wire_switch_in_stage7[121]), .inData_122(wire_switch_in_stage7[122]), .inData_123(wire_switch_in_stage7[123]), .inData_124(wire_switch_in_stage7[124]), .inData_125(wire_switch_in_stage7[125]), .inData_126(wire_switch_in_stage7[126]), .inData_127(wire_switch_in_stage7[127]), .inData_128(wire_switch_in_stage7[128]), .inData_129(wire_switch_in_stage7[129]), .inData_130(wire_switch_in_stage7[130]), .inData_131(wire_switch_in_stage7[131]), .inData_132(wire_switch_in_stage7[132]), .inData_133(wire_switch_in_stage7[133]), .inData_134(wire_switch_in_stage7[134]), .inData_135(wire_switch_in_stage7[135]), .inData_136(wire_switch_in_stage7[136]), .inData_137(wire_switch_in_stage7[137]), .inData_138(wire_switch_in_stage7[138]), .inData_139(wire_switch_in_stage7[139]), .inData_140(wire_switch_in_stage7[140]), .inData_141(wire_switch_in_stage7[141]), .inData_142(wire_switch_in_stage7[142]), .inData_143(wire_switch_in_stage7[143]), .inData_144(wire_switch_in_stage7[144]), .inData_145(wire_switch_in_stage7[145]), .inData_146(wire_switch_in_stage7[146]), .inData_147(wire_switch_in_stage7[147]), .inData_148(wire_switch_in_stage7[148]), .inData_149(wire_switch_in_stage7[149]), .inData_150(wire_switch_in_stage7[150]), .inData_151(wire_switch_in_stage7[151]), .inData_152(wire_switch_in_stage7[152]), .inData_153(wire_switch_in_stage7[153]), .inData_154(wire_switch_in_stage7[154]), .inData_155(wire_switch_in_stage7[155]), .inData_156(wire_switch_in_stage7[156]), .inData_157(wire_switch_in_stage7[157]), .inData_158(wire_switch_in_stage7[158]), .inData_159(wire_switch_in_stage7[159]), .inData_160(wire_switch_in_stage7[160]), .inData_161(wire_switch_in_stage7[161]), .inData_162(wire_switch_in_stage7[162]), .inData_163(wire_switch_in_stage7[163]), .inData_164(wire_switch_in_stage7[164]), .inData_165(wire_switch_in_stage7[165]), .inData_166(wire_switch_in_stage7[166]), .inData_167(wire_switch_in_stage7[167]), .inData_168(wire_switch_in_stage7[168]), .inData_169(wire_switch_in_stage7[169]), .inData_170(wire_switch_in_stage7[170]), .inData_171(wire_switch_in_stage7[171]), .inData_172(wire_switch_in_stage7[172]), .inData_173(wire_switch_in_stage7[173]), .inData_174(wire_switch_in_stage7[174]), .inData_175(wire_switch_in_stage7[175]), .inData_176(wire_switch_in_stage7[176]), .inData_177(wire_switch_in_stage7[177]), .inData_178(wire_switch_in_stage7[178]), .inData_179(wire_switch_in_stage7[179]), .inData_180(wire_switch_in_stage7[180]), .inData_181(wire_switch_in_stage7[181]), .inData_182(wire_switch_in_stage7[182]), .inData_183(wire_switch_in_stage7[183]), .inData_184(wire_switch_in_stage7[184]), .inData_185(wire_switch_in_stage7[185]), .inData_186(wire_switch_in_stage7[186]), .inData_187(wire_switch_in_stage7[187]), .inData_188(wire_switch_in_stage7[188]), .inData_189(wire_switch_in_stage7[189]), .inData_190(wire_switch_in_stage7[190]), .inData_191(wire_switch_in_stage7[191]), .inData_192(wire_switch_in_stage7[192]), .inData_193(wire_switch_in_stage7[193]), .inData_194(wire_switch_in_stage7[194]), .inData_195(wire_switch_in_stage7[195]), .inData_196(wire_switch_in_stage7[196]), .inData_197(wire_switch_in_stage7[197]), .inData_198(wire_switch_in_stage7[198]), .inData_199(wire_switch_in_stage7[199]), .inData_200(wire_switch_in_stage7[200]), .inData_201(wire_switch_in_stage7[201]), .inData_202(wire_switch_in_stage7[202]), .inData_203(wire_switch_in_stage7[203]), .inData_204(wire_switch_in_stage7[204]), .inData_205(wire_switch_in_stage7[205]), .inData_206(wire_switch_in_stage7[206]), .inData_207(wire_switch_in_stage7[207]), .inData_208(wire_switch_in_stage7[208]), .inData_209(wire_switch_in_stage7[209]), .inData_210(wire_switch_in_stage7[210]), .inData_211(wire_switch_in_stage7[211]), .inData_212(wire_switch_in_stage7[212]), .inData_213(wire_switch_in_stage7[213]), .inData_214(wire_switch_in_stage7[214]), .inData_215(wire_switch_in_stage7[215]), .inData_216(wire_switch_in_stage7[216]), .inData_217(wire_switch_in_stage7[217]), .inData_218(wire_switch_in_stage7[218]), .inData_219(wire_switch_in_stage7[219]), .inData_220(wire_switch_in_stage7[220]), .inData_221(wire_switch_in_stage7[221]), .inData_222(wire_switch_in_stage7[222]), .inData_223(wire_switch_in_stage7[223]), .inData_224(wire_switch_in_stage7[224]), .inData_225(wire_switch_in_stage7[225]), .inData_226(wire_switch_in_stage7[226]), .inData_227(wire_switch_in_stage7[227]), .inData_228(wire_switch_in_stage7[228]), .inData_229(wire_switch_in_stage7[229]), .inData_230(wire_switch_in_stage7[230]), .inData_231(wire_switch_in_stage7[231]), .inData_232(wire_switch_in_stage7[232]), .inData_233(wire_switch_in_stage7[233]), .inData_234(wire_switch_in_stage7[234]), .inData_235(wire_switch_in_stage7[235]), .inData_236(wire_switch_in_stage7[236]), .inData_237(wire_switch_in_stage7[237]), .inData_238(wire_switch_in_stage7[238]), .inData_239(wire_switch_in_stage7[239]), .inData_240(wire_switch_in_stage7[240]), .inData_241(wire_switch_in_stage7[241]), .inData_242(wire_switch_in_stage7[242]), .inData_243(wire_switch_in_stage7[243]), .inData_244(wire_switch_in_stage7[244]), .inData_245(wire_switch_in_stage7[245]), .inData_246(wire_switch_in_stage7[246]), .inData_247(wire_switch_in_stage7[247]), .inData_248(wire_switch_in_stage7[248]), .inData_249(wire_switch_in_stage7[249]), .inData_250(wire_switch_in_stage7[250]), .inData_251(wire_switch_in_stage7[251]), .inData_252(wire_switch_in_stage7[252]), .inData_253(wire_switch_in_stage7[253]), .inData_254(wire_switch_in_stage7[254]), .inData_255(wire_switch_in_stage7[255]), 
        .outData_0(wire_switch_out_stage7[0]), .outData_1(wire_switch_out_stage7[1]), .outData_2(wire_switch_out_stage7[2]), .outData_3(wire_switch_out_stage7[3]), .outData_4(wire_switch_out_stage7[4]), .outData_5(wire_switch_out_stage7[5]), .outData_6(wire_switch_out_stage7[6]), .outData_7(wire_switch_out_stage7[7]), .outData_8(wire_switch_out_stage7[8]), .outData_9(wire_switch_out_stage7[9]), .outData_10(wire_switch_out_stage7[10]), .outData_11(wire_switch_out_stage7[11]), .outData_12(wire_switch_out_stage7[12]), .outData_13(wire_switch_out_stage7[13]), .outData_14(wire_switch_out_stage7[14]), .outData_15(wire_switch_out_stage7[15]), .outData_16(wire_switch_out_stage7[16]), .outData_17(wire_switch_out_stage7[17]), .outData_18(wire_switch_out_stage7[18]), .outData_19(wire_switch_out_stage7[19]), .outData_20(wire_switch_out_stage7[20]), .outData_21(wire_switch_out_stage7[21]), .outData_22(wire_switch_out_stage7[22]), .outData_23(wire_switch_out_stage7[23]), .outData_24(wire_switch_out_stage7[24]), .outData_25(wire_switch_out_stage7[25]), .outData_26(wire_switch_out_stage7[26]), .outData_27(wire_switch_out_stage7[27]), .outData_28(wire_switch_out_stage7[28]), .outData_29(wire_switch_out_stage7[29]), .outData_30(wire_switch_out_stage7[30]), .outData_31(wire_switch_out_stage7[31]), .outData_32(wire_switch_out_stage7[32]), .outData_33(wire_switch_out_stage7[33]), .outData_34(wire_switch_out_stage7[34]), .outData_35(wire_switch_out_stage7[35]), .outData_36(wire_switch_out_stage7[36]), .outData_37(wire_switch_out_stage7[37]), .outData_38(wire_switch_out_stage7[38]), .outData_39(wire_switch_out_stage7[39]), .outData_40(wire_switch_out_stage7[40]), .outData_41(wire_switch_out_stage7[41]), .outData_42(wire_switch_out_stage7[42]), .outData_43(wire_switch_out_stage7[43]), .outData_44(wire_switch_out_stage7[44]), .outData_45(wire_switch_out_stage7[45]), .outData_46(wire_switch_out_stage7[46]), .outData_47(wire_switch_out_stage7[47]), .outData_48(wire_switch_out_stage7[48]), .outData_49(wire_switch_out_stage7[49]), .outData_50(wire_switch_out_stage7[50]), .outData_51(wire_switch_out_stage7[51]), .outData_52(wire_switch_out_stage7[52]), .outData_53(wire_switch_out_stage7[53]), .outData_54(wire_switch_out_stage7[54]), .outData_55(wire_switch_out_stage7[55]), .outData_56(wire_switch_out_stage7[56]), .outData_57(wire_switch_out_stage7[57]), .outData_58(wire_switch_out_stage7[58]), .outData_59(wire_switch_out_stage7[59]), .outData_60(wire_switch_out_stage7[60]), .outData_61(wire_switch_out_stage7[61]), .outData_62(wire_switch_out_stage7[62]), .outData_63(wire_switch_out_stage7[63]), .outData_64(wire_switch_out_stage7[64]), .outData_65(wire_switch_out_stage7[65]), .outData_66(wire_switch_out_stage7[66]), .outData_67(wire_switch_out_stage7[67]), .outData_68(wire_switch_out_stage7[68]), .outData_69(wire_switch_out_stage7[69]), .outData_70(wire_switch_out_stage7[70]), .outData_71(wire_switch_out_stage7[71]), .outData_72(wire_switch_out_stage7[72]), .outData_73(wire_switch_out_stage7[73]), .outData_74(wire_switch_out_stage7[74]), .outData_75(wire_switch_out_stage7[75]), .outData_76(wire_switch_out_stage7[76]), .outData_77(wire_switch_out_stage7[77]), .outData_78(wire_switch_out_stage7[78]), .outData_79(wire_switch_out_stage7[79]), .outData_80(wire_switch_out_stage7[80]), .outData_81(wire_switch_out_stage7[81]), .outData_82(wire_switch_out_stage7[82]), .outData_83(wire_switch_out_stage7[83]), .outData_84(wire_switch_out_stage7[84]), .outData_85(wire_switch_out_stage7[85]), .outData_86(wire_switch_out_stage7[86]), .outData_87(wire_switch_out_stage7[87]), .outData_88(wire_switch_out_stage7[88]), .outData_89(wire_switch_out_stage7[89]), .outData_90(wire_switch_out_stage7[90]), .outData_91(wire_switch_out_stage7[91]), .outData_92(wire_switch_out_stage7[92]), .outData_93(wire_switch_out_stage7[93]), .outData_94(wire_switch_out_stage7[94]), .outData_95(wire_switch_out_stage7[95]), .outData_96(wire_switch_out_stage7[96]), .outData_97(wire_switch_out_stage7[97]), .outData_98(wire_switch_out_stage7[98]), .outData_99(wire_switch_out_stage7[99]), .outData_100(wire_switch_out_stage7[100]), .outData_101(wire_switch_out_stage7[101]), .outData_102(wire_switch_out_stage7[102]), .outData_103(wire_switch_out_stage7[103]), .outData_104(wire_switch_out_stage7[104]), .outData_105(wire_switch_out_stage7[105]), .outData_106(wire_switch_out_stage7[106]), .outData_107(wire_switch_out_stage7[107]), .outData_108(wire_switch_out_stage7[108]), .outData_109(wire_switch_out_stage7[109]), .outData_110(wire_switch_out_stage7[110]), .outData_111(wire_switch_out_stage7[111]), .outData_112(wire_switch_out_stage7[112]), .outData_113(wire_switch_out_stage7[113]), .outData_114(wire_switch_out_stage7[114]), .outData_115(wire_switch_out_stage7[115]), .outData_116(wire_switch_out_stage7[116]), .outData_117(wire_switch_out_stage7[117]), .outData_118(wire_switch_out_stage7[118]), .outData_119(wire_switch_out_stage7[119]), .outData_120(wire_switch_out_stage7[120]), .outData_121(wire_switch_out_stage7[121]), .outData_122(wire_switch_out_stage7[122]), .outData_123(wire_switch_out_stage7[123]), .outData_124(wire_switch_out_stage7[124]), .outData_125(wire_switch_out_stage7[125]), .outData_126(wire_switch_out_stage7[126]), .outData_127(wire_switch_out_stage7[127]), .outData_128(wire_switch_out_stage7[128]), .outData_129(wire_switch_out_stage7[129]), .outData_130(wire_switch_out_stage7[130]), .outData_131(wire_switch_out_stage7[131]), .outData_132(wire_switch_out_stage7[132]), .outData_133(wire_switch_out_stage7[133]), .outData_134(wire_switch_out_stage7[134]), .outData_135(wire_switch_out_stage7[135]), .outData_136(wire_switch_out_stage7[136]), .outData_137(wire_switch_out_stage7[137]), .outData_138(wire_switch_out_stage7[138]), .outData_139(wire_switch_out_stage7[139]), .outData_140(wire_switch_out_stage7[140]), .outData_141(wire_switch_out_stage7[141]), .outData_142(wire_switch_out_stage7[142]), .outData_143(wire_switch_out_stage7[143]), .outData_144(wire_switch_out_stage7[144]), .outData_145(wire_switch_out_stage7[145]), .outData_146(wire_switch_out_stage7[146]), .outData_147(wire_switch_out_stage7[147]), .outData_148(wire_switch_out_stage7[148]), .outData_149(wire_switch_out_stage7[149]), .outData_150(wire_switch_out_stage7[150]), .outData_151(wire_switch_out_stage7[151]), .outData_152(wire_switch_out_stage7[152]), .outData_153(wire_switch_out_stage7[153]), .outData_154(wire_switch_out_stage7[154]), .outData_155(wire_switch_out_stage7[155]), .outData_156(wire_switch_out_stage7[156]), .outData_157(wire_switch_out_stage7[157]), .outData_158(wire_switch_out_stage7[158]), .outData_159(wire_switch_out_stage7[159]), .outData_160(wire_switch_out_stage7[160]), .outData_161(wire_switch_out_stage7[161]), .outData_162(wire_switch_out_stage7[162]), .outData_163(wire_switch_out_stage7[163]), .outData_164(wire_switch_out_stage7[164]), .outData_165(wire_switch_out_stage7[165]), .outData_166(wire_switch_out_stage7[166]), .outData_167(wire_switch_out_stage7[167]), .outData_168(wire_switch_out_stage7[168]), .outData_169(wire_switch_out_stage7[169]), .outData_170(wire_switch_out_stage7[170]), .outData_171(wire_switch_out_stage7[171]), .outData_172(wire_switch_out_stage7[172]), .outData_173(wire_switch_out_stage7[173]), .outData_174(wire_switch_out_stage7[174]), .outData_175(wire_switch_out_stage7[175]), .outData_176(wire_switch_out_stage7[176]), .outData_177(wire_switch_out_stage7[177]), .outData_178(wire_switch_out_stage7[178]), .outData_179(wire_switch_out_stage7[179]), .outData_180(wire_switch_out_stage7[180]), .outData_181(wire_switch_out_stage7[181]), .outData_182(wire_switch_out_stage7[182]), .outData_183(wire_switch_out_stage7[183]), .outData_184(wire_switch_out_stage7[184]), .outData_185(wire_switch_out_stage7[185]), .outData_186(wire_switch_out_stage7[186]), .outData_187(wire_switch_out_stage7[187]), .outData_188(wire_switch_out_stage7[188]), .outData_189(wire_switch_out_stage7[189]), .outData_190(wire_switch_out_stage7[190]), .outData_191(wire_switch_out_stage7[191]), .outData_192(wire_switch_out_stage7[192]), .outData_193(wire_switch_out_stage7[193]), .outData_194(wire_switch_out_stage7[194]), .outData_195(wire_switch_out_stage7[195]), .outData_196(wire_switch_out_stage7[196]), .outData_197(wire_switch_out_stage7[197]), .outData_198(wire_switch_out_stage7[198]), .outData_199(wire_switch_out_stage7[199]), .outData_200(wire_switch_out_stage7[200]), .outData_201(wire_switch_out_stage7[201]), .outData_202(wire_switch_out_stage7[202]), .outData_203(wire_switch_out_stage7[203]), .outData_204(wire_switch_out_stage7[204]), .outData_205(wire_switch_out_stage7[205]), .outData_206(wire_switch_out_stage7[206]), .outData_207(wire_switch_out_stage7[207]), .outData_208(wire_switch_out_stage7[208]), .outData_209(wire_switch_out_stage7[209]), .outData_210(wire_switch_out_stage7[210]), .outData_211(wire_switch_out_stage7[211]), .outData_212(wire_switch_out_stage7[212]), .outData_213(wire_switch_out_stage7[213]), .outData_214(wire_switch_out_stage7[214]), .outData_215(wire_switch_out_stage7[215]), .outData_216(wire_switch_out_stage7[216]), .outData_217(wire_switch_out_stage7[217]), .outData_218(wire_switch_out_stage7[218]), .outData_219(wire_switch_out_stage7[219]), .outData_220(wire_switch_out_stage7[220]), .outData_221(wire_switch_out_stage7[221]), .outData_222(wire_switch_out_stage7[222]), .outData_223(wire_switch_out_stage7[223]), .outData_224(wire_switch_out_stage7[224]), .outData_225(wire_switch_out_stage7[225]), .outData_226(wire_switch_out_stage7[226]), .outData_227(wire_switch_out_stage7[227]), .outData_228(wire_switch_out_stage7[228]), .outData_229(wire_switch_out_stage7[229]), .outData_230(wire_switch_out_stage7[230]), .outData_231(wire_switch_out_stage7[231]), .outData_232(wire_switch_out_stage7[232]), .outData_233(wire_switch_out_stage7[233]), .outData_234(wire_switch_out_stage7[234]), .outData_235(wire_switch_out_stage7[235]), .outData_236(wire_switch_out_stage7[236]), .outData_237(wire_switch_out_stage7[237]), .outData_238(wire_switch_out_stage7[238]), .outData_239(wire_switch_out_stage7[239]), .outData_240(wire_switch_out_stage7[240]), .outData_241(wire_switch_out_stage7[241]), .outData_242(wire_switch_out_stage7[242]), .outData_243(wire_switch_out_stage7[243]), .outData_244(wire_switch_out_stage7[244]), .outData_245(wire_switch_out_stage7[245]), .outData_246(wire_switch_out_stage7[246]), .outData_247(wire_switch_out_stage7[247]), .outData_248(wire_switch_out_stage7[248]), .outData_249(wire_switch_out_stage7[249]), .outData_250(wire_switch_out_stage7[250]), .outData_251(wire_switch_out_stage7[251]), .outData_252(wire_switch_out_stage7[252]), .outData_253(wire_switch_out_stage7[253]), .outData_254(wire_switch_out_stage7[254]), .outData_255(wire_switch_out_stage7[255]), 
        .in_start(con_in_start_stage7), .out_start(in_start_stage6), .ctrl(wire_ctrl_stage7), .clk(clk), .rst(rst));
  
  wireCon_dp256_st7_R wire_stage_7(
        .inData_0(wireIn[0]), .inData_1(wireIn[1]), .inData_2(wireIn[2]), .inData_3(wireIn[3]), .inData_4(wireIn[4]), .inData_5(wireIn[5]), .inData_6(wireIn[6]), .inData_7(wireIn[7]), .inData_8(wireIn[8]), .inData_9(wireIn[9]), .inData_10(wireIn[10]), .inData_11(wireIn[11]), .inData_12(wireIn[12]), .inData_13(wireIn[13]), .inData_14(wireIn[14]), .inData_15(wireIn[15]), .inData_16(wireIn[16]), .inData_17(wireIn[17]), .inData_18(wireIn[18]), .inData_19(wireIn[19]), .inData_20(wireIn[20]), .inData_21(wireIn[21]), .inData_22(wireIn[22]), .inData_23(wireIn[23]), .inData_24(wireIn[24]), .inData_25(wireIn[25]), .inData_26(wireIn[26]), .inData_27(wireIn[27]), .inData_28(wireIn[28]), .inData_29(wireIn[29]), .inData_30(wireIn[30]), .inData_31(wireIn[31]), .inData_32(wireIn[32]), .inData_33(wireIn[33]), .inData_34(wireIn[34]), .inData_35(wireIn[35]), .inData_36(wireIn[36]), .inData_37(wireIn[37]), .inData_38(wireIn[38]), .inData_39(wireIn[39]), .inData_40(wireIn[40]), .inData_41(wireIn[41]), .inData_42(wireIn[42]), .inData_43(wireIn[43]), .inData_44(wireIn[44]), .inData_45(wireIn[45]), .inData_46(wireIn[46]), .inData_47(wireIn[47]), .inData_48(wireIn[48]), .inData_49(wireIn[49]), .inData_50(wireIn[50]), .inData_51(wireIn[51]), .inData_52(wireIn[52]), .inData_53(wireIn[53]), .inData_54(wireIn[54]), .inData_55(wireIn[55]), .inData_56(wireIn[56]), .inData_57(wireIn[57]), .inData_58(wireIn[58]), .inData_59(wireIn[59]), .inData_60(wireIn[60]), .inData_61(wireIn[61]), .inData_62(wireIn[62]), .inData_63(wireIn[63]), .inData_64(wireIn[64]), .inData_65(wireIn[65]), .inData_66(wireIn[66]), .inData_67(wireIn[67]), .inData_68(wireIn[68]), .inData_69(wireIn[69]), .inData_70(wireIn[70]), .inData_71(wireIn[71]), .inData_72(wireIn[72]), .inData_73(wireIn[73]), .inData_74(wireIn[74]), .inData_75(wireIn[75]), .inData_76(wireIn[76]), .inData_77(wireIn[77]), .inData_78(wireIn[78]), .inData_79(wireIn[79]), .inData_80(wireIn[80]), .inData_81(wireIn[81]), .inData_82(wireIn[82]), .inData_83(wireIn[83]), .inData_84(wireIn[84]), .inData_85(wireIn[85]), .inData_86(wireIn[86]), .inData_87(wireIn[87]), .inData_88(wireIn[88]), .inData_89(wireIn[89]), .inData_90(wireIn[90]), .inData_91(wireIn[91]), .inData_92(wireIn[92]), .inData_93(wireIn[93]), .inData_94(wireIn[94]), .inData_95(wireIn[95]), .inData_96(wireIn[96]), .inData_97(wireIn[97]), .inData_98(wireIn[98]), .inData_99(wireIn[99]), .inData_100(wireIn[100]), .inData_101(wireIn[101]), .inData_102(wireIn[102]), .inData_103(wireIn[103]), .inData_104(wireIn[104]), .inData_105(wireIn[105]), .inData_106(wireIn[106]), .inData_107(wireIn[107]), .inData_108(wireIn[108]), .inData_109(wireIn[109]), .inData_110(wireIn[110]), .inData_111(wireIn[111]), .inData_112(wireIn[112]), .inData_113(wireIn[113]), .inData_114(wireIn[114]), .inData_115(wireIn[115]), .inData_116(wireIn[116]), .inData_117(wireIn[117]), .inData_118(wireIn[118]), .inData_119(wireIn[119]), .inData_120(wireIn[120]), .inData_121(wireIn[121]), .inData_122(wireIn[122]), .inData_123(wireIn[123]), .inData_124(wireIn[124]), .inData_125(wireIn[125]), .inData_126(wireIn[126]), .inData_127(wireIn[127]), .inData_128(wireIn[128]), .inData_129(wireIn[129]), .inData_130(wireIn[130]), .inData_131(wireIn[131]), .inData_132(wireIn[132]), .inData_133(wireIn[133]), .inData_134(wireIn[134]), .inData_135(wireIn[135]), .inData_136(wireIn[136]), .inData_137(wireIn[137]), .inData_138(wireIn[138]), .inData_139(wireIn[139]), .inData_140(wireIn[140]), .inData_141(wireIn[141]), .inData_142(wireIn[142]), .inData_143(wireIn[143]), .inData_144(wireIn[144]), .inData_145(wireIn[145]), .inData_146(wireIn[146]), .inData_147(wireIn[147]), .inData_148(wireIn[148]), .inData_149(wireIn[149]), .inData_150(wireIn[150]), .inData_151(wireIn[151]), .inData_152(wireIn[152]), .inData_153(wireIn[153]), .inData_154(wireIn[154]), .inData_155(wireIn[155]), .inData_156(wireIn[156]), .inData_157(wireIn[157]), .inData_158(wireIn[158]), .inData_159(wireIn[159]), .inData_160(wireIn[160]), .inData_161(wireIn[161]), .inData_162(wireIn[162]), .inData_163(wireIn[163]), .inData_164(wireIn[164]), .inData_165(wireIn[165]), .inData_166(wireIn[166]), .inData_167(wireIn[167]), .inData_168(wireIn[168]), .inData_169(wireIn[169]), .inData_170(wireIn[170]), .inData_171(wireIn[171]), .inData_172(wireIn[172]), .inData_173(wireIn[173]), .inData_174(wireIn[174]), .inData_175(wireIn[175]), .inData_176(wireIn[176]), .inData_177(wireIn[177]), .inData_178(wireIn[178]), .inData_179(wireIn[179]), .inData_180(wireIn[180]), .inData_181(wireIn[181]), .inData_182(wireIn[182]), .inData_183(wireIn[183]), .inData_184(wireIn[184]), .inData_185(wireIn[185]), .inData_186(wireIn[186]), .inData_187(wireIn[187]), .inData_188(wireIn[188]), .inData_189(wireIn[189]), .inData_190(wireIn[190]), .inData_191(wireIn[191]), .inData_192(wireIn[192]), .inData_193(wireIn[193]), .inData_194(wireIn[194]), .inData_195(wireIn[195]), .inData_196(wireIn[196]), .inData_197(wireIn[197]), .inData_198(wireIn[198]), .inData_199(wireIn[199]), .inData_200(wireIn[200]), .inData_201(wireIn[201]), .inData_202(wireIn[202]), .inData_203(wireIn[203]), .inData_204(wireIn[204]), .inData_205(wireIn[205]), .inData_206(wireIn[206]), .inData_207(wireIn[207]), .inData_208(wireIn[208]), .inData_209(wireIn[209]), .inData_210(wireIn[210]), .inData_211(wireIn[211]), .inData_212(wireIn[212]), .inData_213(wireIn[213]), .inData_214(wireIn[214]), .inData_215(wireIn[215]), .inData_216(wireIn[216]), .inData_217(wireIn[217]), .inData_218(wireIn[218]), .inData_219(wireIn[219]), .inData_220(wireIn[220]), .inData_221(wireIn[221]), .inData_222(wireIn[222]), .inData_223(wireIn[223]), .inData_224(wireIn[224]), .inData_225(wireIn[225]), .inData_226(wireIn[226]), .inData_227(wireIn[227]), .inData_228(wireIn[228]), .inData_229(wireIn[229]), .inData_230(wireIn[230]), .inData_231(wireIn[231]), .inData_232(wireIn[232]), .inData_233(wireIn[233]), .inData_234(wireIn[234]), .inData_235(wireIn[235]), .inData_236(wireIn[236]), .inData_237(wireIn[237]), .inData_238(wireIn[238]), .inData_239(wireIn[239]), .inData_240(wireIn[240]), .inData_241(wireIn[241]), .inData_242(wireIn[242]), .inData_243(wireIn[243]), .inData_244(wireIn[244]), .inData_245(wireIn[245]), .inData_246(wireIn[246]), .inData_247(wireIn[247]), .inData_248(wireIn[248]), .inData_249(wireIn[249]), .inData_250(wireIn[250]), .inData_251(wireIn[251]), .inData_252(wireIn[252]), .inData_253(wireIn[253]), .inData_254(wireIn[254]), .inData_255(wireIn[255]), 
        .outData_0(wire_switch_in_stage7[0]), .outData_1(wire_switch_in_stage7[1]), .outData_2(wire_switch_in_stage7[2]), .outData_3(wire_switch_in_stage7[3]), .outData_4(wire_switch_in_stage7[4]), .outData_5(wire_switch_in_stage7[5]), .outData_6(wire_switch_in_stage7[6]), .outData_7(wire_switch_in_stage7[7]), .outData_8(wire_switch_in_stage7[8]), .outData_9(wire_switch_in_stage7[9]), .outData_10(wire_switch_in_stage7[10]), .outData_11(wire_switch_in_stage7[11]), .outData_12(wire_switch_in_stage7[12]), .outData_13(wire_switch_in_stage7[13]), .outData_14(wire_switch_in_stage7[14]), .outData_15(wire_switch_in_stage7[15]), .outData_16(wire_switch_in_stage7[16]), .outData_17(wire_switch_in_stage7[17]), .outData_18(wire_switch_in_stage7[18]), .outData_19(wire_switch_in_stage7[19]), .outData_20(wire_switch_in_stage7[20]), .outData_21(wire_switch_in_stage7[21]), .outData_22(wire_switch_in_stage7[22]), .outData_23(wire_switch_in_stage7[23]), .outData_24(wire_switch_in_stage7[24]), .outData_25(wire_switch_in_stage7[25]), .outData_26(wire_switch_in_stage7[26]), .outData_27(wire_switch_in_stage7[27]), .outData_28(wire_switch_in_stage7[28]), .outData_29(wire_switch_in_stage7[29]), .outData_30(wire_switch_in_stage7[30]), .outData_31(wire_switch_in_stage7[31]), .outData_32(wire_switch_in_stage7[32]), .outData_33(wire_switch_in_stage7[33]), .outData_34(wire_switch_in_stage7[34]), .outData_35(wire_switch_in_stage7[35]), .outData_36(wire_switch_in_stage7[36]), .outData_37(wire_switch_in_stage7[37]), .outData_38(wire_switch_in_stage7[38]), .outData_39(wire_switch_in_stage7[39]), .outData_40(wire_switch_in_stage7[40]), .outData_41(wire_switch_in_stage7[41]), .outData_42(wire_switch_in_stage7[42]), .outData_43(wire_switch_in_stage7[43]), .outData_44(wire_switch_in_stage7[44]), .outData_45(wire_switch_in_stage7[45]), .outData_46(wire_switch_in_stage7[46]), .outData_47(wire_switch_in_stage7[47]), .outData_48(wire_switch_in_stage7[48]), .outData_49(wire_switch_in_stage7[49]), .outData_50(wire_switch_in_stage7[50]), .outData_51(wire_switch_in_stage7[51]), .outData_52(wire_switch_in_stage7[52]), .outData_53(wire_switch_in_stage7[53]), .outData_54(wire_switch_in_stage7[54]), .outData_55(wire_switch_in_stage7[55]), .outData_56(wire_switch_in_stage7[56]), .outData_57(wire_switch_in_stage7[57]), .outData_58(wire_switch_in_stage7[58]), .outData_59(wire_switch_in_stage7[59]), .outData_60(wire_switch_in_stage7[60]), .outData_61(wire_switch_in_stage7[61]), .outData_62(wire_switch_in_stage7[62]), .outData_63(wire_switch_in_stage7[63]), .outData_64(wire_switch_in_stage7[64]), .outData_65(wire_switch_in_stage7[65]), .outData_66(wire_switch_in_stage7[66]), .outData_67(wire_switch_in_stage7[67]), .outData_68(wire_switch_in_stage7[68]), .outData_69(wire_switch_in_stage7[69]), .outData_70(wire_switch_in_stage7[70]), .outData_71(wire_switch_in_stage7[71]), .outData_72(wire_switch_in_stage7[72]), .outData_73(wire_switch_in_stage7[73]), .outData_74(wire_switch_in_stage7[74]), .outData_75(wire_switch_in_stage7[75]), .outData_76(wire_switch_in_stage7[76]), .outData_77(wire_switch_in_stage7[77]), .outData_78(wire_switch_in_stage7[78]), .outData_79(wire_switch_in_stage7[79]), .outData_80(wire_switch_in_stage7[80]), .outData_81(wire_switch_in_stage7[81]), .outData_82(wire_switch_in_stage7[82]), .outData_83(wire_switch_in_stage7[83]), .outData_84(wire_switch_in_stage7[84]), .outData_85(wire_switch_in_stage7[85]), .outData_86(wire_switch_in_stage7[86]), .outData_87(wire_switch_in_stage7[87]), .outData_88(wire_switch_in_stage7[88]), .outData_89(wire_switch_in_stage7[89]), .outData_90(wire_switch_in_stage7[90]), .outData_91(wire_switch_in_stage7[91]), .outData_92(wire_switch_in_stage7[92]), .outData_93(wire_switch_in_stage7[93]), .outData_94(wire_switch_in_stage7[94]), .outData_95(wire_switch_in_stage7[95]), .outData_96(wire_switch_in_stage7[96]), .outData_97(wire_switch_in_stage7[97]), .outData_98(wire_switch_in_stage7[98]), .outData_99(wire_switch_in_stage7[99]), .outData_100(wire_switch_in_stage7[100]), .outData_101(wire_switch_in_stage7[101]), .outData_102(wire_switch_in_stage7[102]), .outData_103(wire_switch_in_stage7[103]), .outData_104(wire_switch_in_stage7[104]), .outData_105(wire_switch_in_stage7[105]), .outData_106(wire_switch_in_stage7[106]), .outData_107(wire_switch_in_stage7[107]), .outData_108(wire_switch_in_stage7[108]), .outData_109(wire_switch_in_stage7[109]), .outData_110(wire_switch_in_stage7[110]), .outData_111(wire_switch_in_stage7[111]), .outData_112(wire_switch_in_stage7[112]), .outData_113(wire_switch_in_stage7[113]), .outData_114(wire_switch_in_stage7[114]), .outData_115(wire_switch_in_stage7[115]), .outData_116(wire_switch_in_stage7[116]), .outData_117(wire_switch_in_stage7[117]), .outData_118(wire_switch_in_stage7[118]), .outData_119(wire_switch_in_stage7[119]), .outData_120(wire_switch_in_stage7[120]), .outData_121(wire_switch_in_stage7[121]), .outData_122(wire_switch_in_stage7[122]), .outData_123(wire_switch_in_stage7[123]), .outData_124(wire_switch_in_stage7[124]), .outData_125(wire_switch_in_stage7[125]), .outData_126(wire_switch_in_stage7[126]), .outData_127(wire_switch_in_stage7[127]), .outData_128(wire_switch_in_stage7[128]), .outData_129(wire_switch_in_stage7[129]), .outData_130(wire_switch_in_stage7[130]), .outData_131(wire_switch_in_stage7[131]), .outData_132(wire_switch_in_stage7[132]), .outData_133(wire_switch_in_stage7[133]), .outData_134(wire_switch_in_stage7[134]), .outData_135(wire_switch_in_stage7[135]), .outData_136(wire_switch_in_stage7[136]), .outData_137(wire_switch_in_stage7[137]), .outData_138(wire_switch_in_stage7[138]), .outData_139(wire_switch_in_stage7[139]), .outData_140(wire_switch_in_stage7[140]), .outData_141(wire_switch_in_stage7[141]), .outData_142(wire_switch_in_stage7[142]), .outData_143(wire_switch_in_stage7[143]), .outData_144(wire_switch_in_stage7[144]), .outData_145(wire_switch_in_stage7[145]), .outData_146(wire_switch_in_stage7[146]), .outData_147(wire_switch_in_stage7[147]), .outData_148(wire_switch_in_stage7[148]), .outData_149(wire_switch_in_stage7[149]), .outData_150(wire_switch_in_stage7[150]), .outData_151(wire_switch_in_stage7[151]), .outData_152(wire_switch_in_stage7[152]), .outData_153(wire_switch_in_stage7[153]), .outData_154(wire_switch_in_stage7[154]), .outData_155(wire_switch_in_stage7[155]), .outData_156(wire_switch_in_stage7[156]), .outData_157(wire_switch_in_stage7[157]), .outData_158(wire_switch_in_stage7[158]), .outData_159(wire_switch_in_stage7[159]), .outData_160(wire_switch_in_stage7[160]), .outData_161(wire_switch_in_stage7[161]), .outData_162(wire_switch_in_stage7[162]), .outData_163(wire_switch_in_stage7[163]), .outData_164(wire_switch_in_stage7[164]), .outData_165(wire_switch_in_stage7[165]), .outData_166(wire_switch_in_stage7[166]), .outData_167(wire_switch_in_stage7[167]), .outData_168(wire_switch_in_stage7[168]), .outData_169(wire_switch_in_stage7[169]), .outData_170(wire_switch_in_stage7[170]), .outData_171(wire_switch_in_stage7[171]), .outData_172(wire_switch_in_stage7[172]), .outData_173(wire_switch_in_stage7[173]), .outData_174(wire_switch_in_stage7[174]), .outData_175(wire_switch_in_stage7[175]), .outData_176(wire_switch_in_stage7[176]), .outData_177(wire_switch_in_stage7[177]), .outData_178(wire_switch_in_stage7[178]), .outData_179(wire_switch_in_stage7[179]), .outData_180(wire_switch_in_stage7[180]), .outData_181(wire_switch_in_stage7[181]), .outData_182(wire_switch_in_stage7[182]), .outData_183(wire_switch_in_stage7[183]), .outData_184(wire_switch_in_stage7[184]), .outData_185(wire_switch_in_stage7[185]), .outData_186(wire_switch_in_stage7[186]), .outData_187(wire_switch_in_stage7[187]), .outData_188(wire_switch_in_stage7[188]), .outData_189(wire_switch_in_stage7[189]), .outData_190(wire_switch_in_stage7[190]), .outData_191(wire_switch_in_stage7[191]), .outData_192(wire_switch_in_stage7[192]), .outData_193(wire_switch_in_stage7[193]), .outData_194(wire_switch_in_stage7[194]), .outData_195(wire_switch_in_stage7[195]), .outData_196(wire_switch_in_stage7[196]), .outData_197(wire_switch_in_stage7[197]), .outData_198(wire_switch_in_stage7[198]), .outData_199(wire_switch_in_stage7[199]), .outData_200(wire_switch_in_stage7[200]), .outData_201(wire_switch_in_stage7[201]), .outData_202(wire_switch_in_stage7[202]), .outData_203(wire_switch_in_stage7[203]), .outData_204(wire_switch_in_stage7[204]), .outData_205(wire_switch_in_stage7[205]), .outData_206(wire_switch_in_stage7[206]), .outData_207(wire_switch_in_stage7[207]), .outData_208(wire_switch_in_stage7[208]), .outData_209(wire_switch_in_stage7[209]), .outData_210(wire_switch_in_stage7[210]), .outData_211(wire_switch_in_stage7[211]), .outData_212(wire_switch_in_stage7[212]), .outData_213(wire_switch_in_stage7[213]), .outData_214(wire_switch_in_stage7[214]), .outData_215(wire_switch_in_stage7[215]), .outData_216(wire_switch_in_stage7[216]), .outData_217(wire_switch_in_stage7[217]), .outData_218(wire_switch_in_stage7[218]), .outData_219(wire_switch_in_stage7[219]), .outData_220(wire_switch_in_stage7[220]), .outData_221(wire_switch_in_stage7[221]), .outData_222(wire_switch_in_stage7[222]), .outData_223(wire_switch_in_stage7[223]), .outData_224(wire_switch_in_stage7[224]), .outData_225(wire_switch_in_stage7[225]), .outData_226(wire_switch_in_stage7[226]), .outData_227(wire_switch_in_stage7[227]), .outData_228(wire_switch_in_stage7[228]), .outData_229(wire_switch_in_stage7[229]), .outData_230(wire_switch_in_stage7[230]), .outData_231(wire_switch_in_stage7[231]), .outData_232(wire_switch_in_stage7[232]), .outData_233(wire_switch_in_stage7[233]), .outData_234(wire_switch_in_stage7[234]), .outData_235(wire_switch_in_stage7[235]), .outData_236(wire_switch_in_stage7[236]), .outData_237(wire_switch_in_stage7[237]), .outData_238(wire_switch_in_stage7[238]), .outData_239(wire_switch_in_stage7[239]), .outData_240(wire_switch_in_stage7[240]), .outData_241(wire_switch_in_stage7[241]), .outData_242(wire_switch_in_stage7[242]), .outData_243(wire_switch_in_stage7[243]), .outData_244(wire_switch_in_stage7[244]), .outData_245(wire_switch_in_stage7[245]), .outData_246(wire_switch_in_stage7[246]), .outData_247(wire_switch_in_stage7[247]), .outData_248(wire_switch_in_stage7[248]), .outData_249(wire_switch_in_stage7[249]), .outData_250(wire_switch_in_stage7[250]), .outData_251(wire_switch_in_stage7[251]), .outData_252(wire_switch_in_stage7[252]), .outData_253(wire_switch_in_stage7[253]), .outData_254(wire_switch_in_stage7[254]), .outData_255(wire_switch_in_stage7[255]), 
        .in_start(in_start_stage7), .out_start(con_in_start_stage7), .clk(clk), .rst(rst)); 

  
  wire [7:0] counter_w;
  assign counter_w = counter_in; 
  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[0] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[1] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[2] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[3] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[4] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[5] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[6] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[7] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[8] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[9] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[10] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[11] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[12] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[13] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[14] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[15] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[16] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[17] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[18] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[19] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[20] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[21] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[22] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[23] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[24] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[25] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[26] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[27] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[28] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[29] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[30] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[31] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[32] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[33] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[34] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[35] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[36] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[37] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[38] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[39] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[40] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[41] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[42] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[43] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[44] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[45] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[46] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[47] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[48] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[49] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[50] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[51] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[52] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[53] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[54] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[55] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[56] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[57] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[58] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[59] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[60] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[61] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[62] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[63] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[64] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[65] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[66] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[67] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[68] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[69] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[70] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[71] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[72] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[73] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[74] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[75] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[76] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[77] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[78] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[79] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[80] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[81] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[82] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[83] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[84] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[85] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[86] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[87] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[88] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[89] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[90] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[91] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[92] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[93] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[94] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[95] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[96] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[97] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[98] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[99] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[100] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[101] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[102] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[103] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[104] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[105] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[106] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[107] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[108] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[109] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[110] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[111] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[112] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[113] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[114] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[115] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[116] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[117] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[118] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[119] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[120] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[121] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[122] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[123] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[124] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[125] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[126] <= counter_w[0]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage7[127] <= counter_w[0]; 
  end                            

  wire [DATA_WIDTH-1:0] wire_switch_in_stage6[255:0];
  wire [DATA_WIDTH-1:0] wire_switch_out_stage6[255:0];
  reg [127:0] wire_ctrl_stage6;

  switches_stage_st6_0_R switch_stage_6(
        .inData_0(wire_switch_in_stage6[0]), .inData_1(wire_switch_in_stage6[1]), .inData_2(wire_switch_in_stage6[2]), .inData_3(wire_switch_in_stage6[3]), .inData_4(wire_switch_in_stage6[4]), .inData_5(wire_switch_in_stage6[5]), .inData_6(wire_switch_in_stage6[6]), .inData_7(wire_switch_in_stage6[7]), .inData_8(wire_switch_in_stage6[8]), .inData_9(wire_switch_in_stage6[9]), .inData_10(wire_switch_in_stage6[10]), .inData_11(wire_switch_in_stage6[11]), .inData_12(wire_switch_in_stage6[12]), .inData_13(wire_switch_in_stage6[13]), .inData_14(wire_switch_in_stage6[14]), .inData_15(wire_switch_in_stage6[15]), .inData_16(wire_switch_in_stage6[16]), .inData_17(wire_switch_in_stage6[17]), .inData_18(wire_switch_in_stage6[18]), .inData_19(wire_switch_in_stage6[19]), .inData_20(wire_switch_in_stage6[20]), .inData_21(wire_switch_in_stage6[21]), .inData_22(wire_switch_in_stage6[22]), .inData_23(wire_switch_in_stage6[23]), .inData_24(wire_switch_in_stage6[24]), .inData_25(wire_switch_in_stage6[25]), .inData_26(wire_switch_in_stage6[26]), .inData_27(wire_switch_in_stage6[27]), .inData_28(wire_switch_in_stage6[28]), .inData_29(wire_switch_in_stage6[29]), .inData_30(wire_switch_in_stage6[30]), .inData_31(wire_switch_in_stage6[31]), .inData_32(wire_switch_in_stage6[32]), .inData_33(wire_switch_in_stage6[33]), .inData_34(wire_switch_in_stage6[34]), .inData_35(wire_switch_in_stage6[35]), .inData_36(wire_switch_in_stage6[36]), .inData_37(wire_switch_in_stage6[37]), .inData_38(wire_switch_in_stage6[38]), .inData_39(wire_switch_in_stage6[39]), .inData_40(wire_switch_in_stage6[40]), .inData_41(wire_switch_in_stage6[41]), .inData_42(wire_switch_in_stage6[42]), .inData_43(wire_switch_in_stage6[43]), .inData_44(wire_switch_in_stage6[44]), .inData_45(wire_switch_in_stage6[45]), .inData_46(wire_switch_in_stage6[46]), .inData_47(wire_switch_in_stage6[47]), .inData_48(wire_switch_in_stage6[48]), .inData_49(wire_switch_in_stage6[49]), .inData_50(wire_switch_in_stage6[50]), .inData_51(wire_switch_in_stage6[51]), .inData_52(wire_switch_in_stage6[52]), .inData_53(wire_switch_in_stage6[53]), .inData_54(wire_switch_in_stage6[54]), .inData_55(wire_switch_in_stage6[55]), .inData_56(wire_switch_in_stage6[56]), .inData_57(wire_switch_in_stage6[57]), .inData_58(wire_switch_in_stage6[58]), .inData_59(wire_switch_in_stage6[59]), .inData_60(wire_switch_in_stage6[60]), .inData_61(wire_switch_in_stage6[61]), .inData_62(wire_switch_in_stage6[62]), .inData_63(wire_switch_in_stage6[63]), .inData_64(wire_switch_in_stage6[64]), .inData_65(wire_switch_in_stage6[65]), .inData_66(wire_switch_in_stage6[66]), .inData_67(wire_switch_in_stage6[67]), .inData_68(wire_switch_in_stage6[68]), .inData_69(wire_switch_in_stage6[69]), .inData_70(wire_switch_in_stage6[70]), .inData_71(wire_switch_in_stage6[71]), .inData_72(wire_switch_in_stage6[72]), .inData_73(wire_switch_in_stage6[73]), .inData_74(wire_switch_in_stage6[74]), .inData_75(wire_switch_in_stage6[75]), .inData_76(wire_switch_in_stage6[76]), .inData_77(wire_switch_in_stage6[77]), .inData_78(wire_switch_in_stage6[78]), .inData_79(wire_switch_in_stage6[79]), .inData_80(wire_switch_in_stage6[80]), .inData_81(wire_switch_in_stage6[81]), .inData_82(wire_switch_in_stage6[82]), .inData_83(wire_switch_in_stage6[83]), .inData_84(wire_switch_in_stage6[84]), .inData_85(wire_switch_in_stage6[85]), .inData_86(wire_switch_in_stage6[86]), .inData_87(wire_switch_in_stage6[87]), .inData_88(wire_switch_in_stage6[88]), .inData_89(wire_switch_in_stage6[89]), .inData_90(wire_switch_in_stage6[90]), .inData_91(wire_switch_in_stage6[91]), .inData_92(wire_switch_in_stage6[92]), .inData_93(wire_switch_in_stage6[93]), .inData_94(wire_switch_in_stage6[94]), .inData_95(wire_switch_in_stage6[95]), .inData_96(wire_switch_in_stage6[96]), .inData_97(wire_switch_in_stage6[97]), .inData_98(wire_switch_in_stage6[98]), .inData_99(wire_switch_in_stage6[99]), .inData_100(wire_switch_in_stage6[100]), .inData_101(wire_switch_in_stage6[101]), .inData_102(wire_switch_in_stage6[102]), .inData_103(wire_switch_in_stage6[103]), .inData_104(wire_switch_in_stage6[104]), .inData_105(wire_switch_in_stage6[105]), .inData_106(wire_switch_in_stage6[106]), .inData_107(wire_switch_in_stage6[107]), .inData_108(wire_switch_in_stage6[108]), .inData_109(wire_switch_in_stage6[109]), .inData_110(wire_switch_in_stage6[110]), .inData_111(wire_switch_in_stage6[111]), .inData_112(wire_switch_in_stage6[112]), .inData_113(wire_switch_in_stage6[113]), .inData_114(wire_switch_in_stage6[114]), .inData_115(wire_switch_in_stage6[115]), .inData_116(wire_switch_in_stage6[116]), .inData_117(wire_switch_in_stage6[117]), .inData_118(wire_switch_in_stage6[118]), .inData_119(wire_switch_in_stage6[119]), .inData_120(wire_switch_in_stage6[120]), .inData_121(wire_switch_in_stage6[121]), .inData_122(wire_switch_in_stage6[122]), .inData_123(wire_switch_in_stage6[123]), .inData_124(wire_switch_in_stage6[124]), .inData_125(wire_switch_in_stage6[125]), .inData_126(wire_switch_in_stage6[126]), .inData_127(wire_switch_in_stage6[127]), .inData_128(wire_switch_in_stage6[128]), .inData_129(wire_switch_in_stage6[129]), .inData_130(wire_switch_in_stage6[130]), .inData_131(wire_switch_in_stage6[131]), .inData_132(wire_switch_in_stage6[132]), .inData_133(wire_switch_in_stage6[133]), .inData_134(wire_switch_in_stage6[134]), .inData_135(wire_switch_in_stage6[135]), .inData_136(wire_switch_in_stage6[136]), .inData_137(wire_switch_in_stage6[137]), .inData_138(wire_switch_in_stage6[138]), .inData_139(wire_switch_in_stage6[139]), .inData_140(wire_switch_in_stage6[140]), .inData_141(wire_switch_in_stage6[141]), .inData_142(wire_switch_in_stage6[142]), .inData_143(wire_switch_in_stage6[143]), .inData_144(wire_switch_in_stage6[144]), .inData_145(wire_switch_in_stage6[145]), .inData_146(wire_switch_in_stage6[146]), .inData_147(wire_switch_in_stage6[147]), .inData_148(wire_switch_in_stage6[148]), .inData_149(wire_switch_in_stage6[149]), .inData_150(wire_switch_in_stage6[150]), .inData_151(wire_switch_in_stage6[151]), .inData_152(wire_switch_in_stage6[152]), .inData_153(wire_switch_in_stage6[153]), .inData_154(wire_switch_in_stage6[154]), .inData_155(wire_switch_in_stage6[155]), .inData_156(wire_switch_in_stage6[156]), .inData_157(wire_switch_in_stage6[157]), .inData_158(wire_switch_in_stage6[158]), .inData_159(wire_switch_in_stage6[159]), .inData_160(wire_switch_in_stage6[160]), .inData_161(wire_switch_in_stage6[161]), .inData_162(wire_switch_in_stage6[162]), .inData_163(wire_switch_in_stage6[163]), .inData_164(wire_switch_in_stage6[164]), .inData_165(wire_switch_in_stage6[165]), .inData_166(wire_switch_in_stage6[166]), .inData_167(wire_switch_in_stage6[167]), .inData_168(wire_switch_in_stage6[168]), .inData_169(wire_switch_in_stage6[169]), .inData_170(wire_switch_in_stage6[170]), .inData_171(wire_switch_in_stage6[171]), .inData_172(wire_switch_in_stage6[172]), .inData_173(wire_switch_in_stage6[173]), .inData_174(wire_switch_in_stage6[174]), .inData_175(wire_switch_in_stage6[175]), .inData_176(wire_switch_in_stage6[176]), .inData_177(wire_switch_in_stage6[177]), .inData_178(wire_switch_in_stage6[178]), .inData_179(wire_switch_in_stage6[179]), .inData_180(wire_switch_in_stage6[180]), .inData_181(wire_switch_in_stage6[181]), .inData_182(wire_switch_in_stage6[182]), .inData_183(wire_switch_in_stage6[183]), .inData_184(wire_switch_in_stage6[184]), .inData_185(wire_switch_in_stage6[185]), .inData_186(wire_switch_in_stage6[186]), .inData_187(wire_switch_in_stage6[187]), .inData_188(wire_switch_in_stage6[188]), .inData_189(wire_switch_in_stage6[189]), .inData_190(wire_switch_in_stage6[190]), .inData_191(wire_switch_in_stage6[191]), .inData_192(wire_switch_in_stage6[192]), .inData_193(wire_switch_in_stage6[193]), .inData_194(wire_switch_in_stage6[194]), .inData_195(wire_switch_in_stage6[195]), .inData_196(wire_switch_in_stage6[196]), .inData_197(wire_switch_in_stage6[197]), .inData_198(wire_switch_in_stage6[198]), .inData_199(wire_switch_in_stage6[199]), .inData_200(wire_switch_in_stage6[200]), .inData_201(wire_switch_in_stage6[201]), .inData_202(wire_switch_in_stage6[202]), .inData_203(wire_switch_in_stage6[203]), .inData_204(wire_switch_in_stage6[204]), .inData_205(wire_switch_in_stage6[205]), .inData_206(wire_switch_in_stage6[206]), .inData_207(wire_switch_in_stage6[207]), .inData_208(wire_switch_in_stage6[208]), .inData_209(wire_switch_in_stage6[209]), .inData_210(wire_switch_in_stage6[210]), .inData_211(wire_switch_in_stage6[211]), .inData_212(wire_switch_in_stage6[212]), .inData_213(wire_switch_in_stage6[213]), .inData_214(wire_switch_in_stage6[214]), .inData_215(wire_switch_in_stage6[215]), .inData_216(wire_switch_in_stage6[216]), .inData_217(wire_switch_in_stage6[217]), .inData_218(wire_switch_in_stage6[218]), .inData_219(wire_switch_in_stage6[219]), .inData_220(wire_switch_in_stage6[220]), .inData_221(wire_switch_in_stage6[221]), .inData_222(wire_switch_in_stage6[222]), .inData_223(wire_switch_in_stage6[223]), .inData_224(wire_switch_in_stage6[224]), .inData_225(wire_switch_in_stage6[225]), .inData_226(wire_switch_in_stage6[226]), .inData_227(wire_switch_in_stage6[227]), .inData_228(wire_switch_in_stage6[228]), .inData_229(wire_switch_in_stage6[229]), .inData_230(wire_switch_in_stage6[230]), .inData_231(wire_switch_in_stage6[231]), .inData_232(wire_switch_in_stage6[232]), .inData_233(wire_switch_in_stage6[233]), .inData_234(wire_switch_in_stage6[234]), .inData_235(wire_switch_in_stage6[235]), .inData_236(wire_switch_in_stage6[236]), .inData_237(wire_switch_in_stage6[237]), .inData_238(wire_switch_in_stage6[238]), .inData_239(wire_switch_in_stage6[239]), .inData_240(wire_switch_in_stage6[240]), .inData_241(wire_switch_in_stage6[241]), .inData_242(wire_switch_in_stage6[242]), .inData_243(wire_switch_in_stage6[243]), .inData_244(wire_switch_in_stage6[244]), .inData_245(wire_switch_in_stage6[245]), .inData_246(wire_switch_in_stage6[246]), .inData_247(wire_switch_in_stage6[247]), .inData_248(wire_switch_in_stage6[248]), .inData_249(wire_switch_in_stage6[249]), .inData_250(wire_switch_in_stage6[250]), .inData_251(wire_switch_in_stage6[251]), .inData_252(wire_switch_in_stage6[252]), .inData_253(wire_switch_in_stage6[253]), .inData_254(wire_switch_in_stage6[254]), .inData_255(wire_switch_in_stage6[255]), 
        .outData_0(wire_switch_out_stage6[0]), .outData_1(wire_switch_out_stage6[1]), .outData_2(wire_switch_out_stage6[2]), .outData_3(wire_switch_out_stage6[3]), .outData_4(wire_switch_out_stage6[4]), .outData_5(wire_switch_out_stage6[5]), .outData_6(wire_switch_out_stage6[6]), .outData_7(wire_switch_out_stage6[7]), .outData_8(wire_switch_out_stage6[8]), .outData_9(wire_switch_out_stage6[9]), .outData_10(wire_switch_out_stage6[10]), .outData_11(wire_switch_out_stage6[11]), .outData_12(wire_switch_out_stage6[12]), .outData_13(wire_switch_out_stage6[13]), .outData_14(wire_switch_out_stage6[14]), .outData_15(wire_switch_out_stage6[15]), .outData_16(wire_switch_out_stage6[16]), .outData_17(wire_switch_out_stage6[17]), .outData_18(wire_switch_out_stage6[18]), .outData_19(wire_switch_out_stage6[19]), .outData_20(wire_switch_out_stage6[20]), .outData_21(wire_switch_out_stage6[21]), .outData_22(wire_switch_out_stage6[22]), .outData_23(wire_switch_out_stage6[23]), .outData_24(wire_switch_out_stage6[24]), .outData_25(wire_switch_out_stage6[25]), .outData_26(wire_switch_out_stage6[26]), .outData_27(wire_switch_out_stage6[27]), .outData_28(wire_switch_out_stage6[28]), .outData_29(wire_switch_out_stage6[29]), .outData_30(wire_switch_out_stage6[30]), .outData_31(wire_switch_out_stage6[31]), .outData_32(wire_switch_out_stage6[32]), .outData_33(wire_switch_out_stage6[33]), .outData_34(wire_switch_out_stage6[34]), .outData_35(wire_switch_out_stage6[35]), .outData_36(wire_switch_out_stage6[36]), .outData_37(wire_switch_out_stage6[37]), .outData_38(wire_switch_out_stage6[38]), .outData_39(wire_switch_out_stage6[39]), .outData_40(wire_switch_out_stage6[40]), .outData_41(wire_switch_out_stage6[41]), .outData_42(wire_switch_out_stage6[42]), .outData_43(wire_switch_out_stage6[43]), .outData_44(wire_switch_out_stage6[44]), .outData_45(wire_switch_out_stage6[45]), .outData_46(wire_switch_out_stage6[46]), .outData_47(wire_switch_out_stage6[47]), .outData_48(wire_switch_out_stage6[48]), .outData_49(wire_switch_out_stage6[49]), .outData_50(wire_switch_out_stage6[50]), .outData_51(wire_switch_out_stage6[51]), .outData_52(wire_switch_out_stage6[52]), .outData_53(wire_switch_out_stage6[53]), .outData_54(wire_switch_out_stage6[54]), .outData_55(wire_switch_out_stage6[55]), .outData_56(wire_switch_out_stage6[56]), .outData_57(wire_switch_out_stage6[57]), .outData_58(wire_switch_out_stage6[58]), .outData_59(wire_switch_out_stage6[59]), .outData_60(wire_switch_out_stage6[60]), .outData_61(wire_switch_out_stage6[61]), .outData_62(wire_switch_out_stage6[62]), .outData_63(wire_switch_out_stage6[63]), .outData_64(wire_switch_out_stage6[64]), .outData_65(wire_switch_out_stage6[65]), .outData_66(wire_switch_out_stage6[66]), .outData_67(wire_switch_out_stage6[67]), .outData_68(wire_switch_out_stage6[68]), .outData_69(wire_switch_out_stage6[69]), .outData_70(wire_switch_out_stage6[70]), .outData_71(wire_switch_out_stage6[71]), .outData_72(wire_switch_out_stage6[72]), .outData_73(wire_switch_out_stage6[73]), .outData_74(wire_switch_out_stage6[74]), .outData_75(wire_switch_out_stage6[75]), .outData_76(wire_switch_out_stage6[76]), .outData_77(wire_switch_out_stage6[77]), .outData_78(wire_switch_out_stage6[78]), .outData_79(wire_switch_out_stage6[79]), .outData_80(wire_switch_out_stage6[80]), .outData_81(wire_switch_out_stage6[81]), .outData_82(wire_switch_out_stage6[82]), .outData_83(wire_switch_out_stage6[83]), .outData_84(wire_switch_out_stage6[84]), .outData_85(wire_switch_out_stage6[85]), .outData_86(wire_switch_out_stage6[86]), .outData_87(wire_switch_out_stage6[87]), .outData_88(wire_switch_out_stage6[88]), .outData_89(wire_switch_out_stage6[89]), .outData_90(wire_switch_out_stage6[90]), .outData_91(wire_switch_out_stage6[91]), .outData_92(wire_switch_out_stage6[92]), .outData_93(wire_switch_out_stage6[93]), .outData_94(wire_switch_out_stage6[94]), .outData_95(wire_switch_out_stage6[95]), .outData_96(wire_switch_out_stage6[96]), .outData_97(wire_switch_out_stage6[97]), .outData_98(wire_switch_out_stage6[98]), .outData_99(wire_switch_out_stage6[99]), .outData_100(wire_switch_out_stage6[100]), .outData_101(wire_switch_out_stage6[101]), .outData_102(wire_switch_out_stage6[102]), .outData_103(wire_switch_out_stage6[103]), .outData_104(wire_switch_out_stage6[104]), .outData_105(wire_switch_out_stage6[105]), .outData_106(wire_switch_out_stage6[106]), .outData_107(wire_switch_out_stage6[107]), .outData_108(wire_switch_out_stage6[108]), .outData_109(wire_switch_out_stage6[109]), .outData_110(wire_switch_out_stage6[110]), .outData_111(wire_switch_out_stage6[111]), .outData_112(wire_switch_out_stage6[112]), .outData_113(wire_switch_out_stage6[113]), .outData_114(wire_switch_out_stage6[114]), .outData_115(wire_switch_out_stage6[115]), .outData_116(wire_switch_out_stage6[116]), .outData_117(wire_switch_out_stage6[117]), .outData_118(wire_switch_out_stage6[118]), .outData_119(wire_switch_out_stage6[119]), .outData_120(wire_switch_out_stage6[120]), .outData_121(wire_switch_out_stage6[121]), .outData_122(wire_switch_out_stage6[122]), .outData_123(wire_switch_out_stage6[123]), .outData_124(wire_switch_out_stage6[124]), .outData_125(wire_switch_out_stage6[125]), .outData_126(wire_switch_out_stage6[126]), .outData_127(wire_switch_out_stage6[127]), .outData_128(wire_switch_out_stage6[128]), .outData_129(wire_switch_out_stage6[129]), .outData_130(wire_switch_out_stage6[130]), .outData_131(wire_switch_out_stage6[131]), .outData_132(wire_switch_out_stage6[132]), .outData_133(wire_switch_out_stage6[133]), .outData_134(wire_switch_out_stage6[134]), .outData_135(wire_switch_out_stage6[135]), .outData_136(wire_switch_out_stage6[136]), .outData_137(wire_switch_out_stage6[137]), .outData_138(wire_switch_out_stage6[138]), .outData_139(wire_switch_out_stage6[139]), .outData_140(wire_switch_out_stage6[140]), .outData_141(wire_switch_out_stage6[141]), .outData_142(wire_switch_out_stage6[142]), .outData_143(wire_switch_out_stage6[143]), .outData_144(wire_switch_out_stage6[144]), .outData_145(wire_switch_out_stage6[145]), .outData_146(wire_switch_out_stage6[146]), .outData_147(wire_switch_out_stage6[147]), .outData_148(wire_switch_out_stage6[148]), .outData_149(wire_switch_out_stage6[149]), .outData_150(wire_switch_out_stage6[150]), .outData_151(wire_switch_out_stage6[151]), .outData_152(wire_switch_out_stage6[152]), .outData_153(wire_switch_out_stage6[153]), .outData_154(wire_switch_out_stage6[154]), .outData_155(wire_switch_out_stage6[155]), .outData_156(wire_switch_out_stage6[156]), .outData_157(wire_switch_out_stage6[157]), .outData_158(wire_switch_out_stage6[158]), .outData_159(wire_switch_out_stage6[159]), .outData_160(wire_switch_out_stage6[160]), .outData_161(wire_switch_out_stage6[161]), .outData_162(wire_switch_out_stage6[162]), .outData_163(wire_switch_out_stage6[163]), .outData_164(wire_switch_out_stage6[164]), .outData_165(wire_switch_out_stage6[165]), .outData_166(wire_switch_out_stage6[166]), .outData_167(wire_switch_out_stage6[167]), .outData_168(wire_switch_out_stage6[168]), .outData_169(wire_switch_out_stage6[169]), .outData_170(wire_switch_out_stage6[170]), .outData_171(wire_switch_out_stage6[171]), .outData_172(wire_switch_out_stage6[172]), .outData_173(wire_switch_out_stage6[173]), .outData_174(wire_switch_out_stage6[174]), .outData_175(wire_switch_out_stage6[175]), .outData_176(wire_switch_out_stage6[176]), .outData_177(wire_switch_out_stage6[177]), .outData_178(wire_switch_out_stage6[178]), .outData_179(wire_switch_out_stage6[179]), .outData_180(wire_switch_out_stage6[180]), .outData_181(wire_switch_out_stage6[181]), .outData_182(wire_switch_out_stage6[182]), .outData_183(wire_switch_out_stage6[183]), .outData_184(wire_switch_out_stage6[184]), .outData_185(wire_switch_out_stage6[185]), .outData_186(wire_switch_out_stage6[186]), .outData_187(wire_switch_out_stage6[187]), .outData_188(wire_switch_out_stage6[188]), .outData_189(wire_switch_out_stage6[189]), .outData_190(wire_switch_out_stage6[190]), .outData_191(wire_switch_out_stage6[191]), .outData_192(wire_switch_out_stage6[192]), .outData_193(wire_switch_out_stage6[193]), .outData_194(wire_switch_out_stage6[194]), .outData_195(wire_switch_out_stage6[195]), .outData_196(wire_switch_out_stage6[196]), .outData_197(wire_switch_out_stage6[197]), .outData_198(wire_switch_out_stage6[198]), .outData_199(wire_switch_out_stage6[199]), .outData_200(wire_switch_out_stage6[200]), .outData_201(wire_switch_out_stage6[201]), .outData_202(wire_switch_out_stage6[202]), .outData_203(wire_switch_out_stage6[203]), .outData_204(wire_switch_out_stage6[204]), .outData_205(wire_switch_out_stage6[205]), .outData_206(wire_switch_out_stage6[206]), .outData_207(wire_switch_out_stage6[207]), .outData_208(wire_switch_out_stage6[208]), .outData_209(wire_switch_out_stage6[209]), .outData_210(wire_switch_out_stage6[210]), .outData_211(wire_switch_out_stage6[211]), .outData_212(wire_switch_out_stage6[212]), .outData_213(wire_switch_out_stage6[213]), .outData_214(wire_switch_out_stage6[214]), .outData_215(wire_switch_out_stage6[215]), .outData_216(wire_switch_out_stage6[216]), .outData_217(wire_switch_out_stage6[217]), .outData_218(wire_switch_out_stage6[218]), .outData_219(wire_switch_out_stage6[219]), .outData_220(wire_switch_out_stage6[220]), .outData_221(wire_switch_out_stage6[221]), .outData_222(wire_switch_out_stage6[222]), .outData_223(wire_switch_out_stage6[223]), .outData_224(wire_switch_out_stage6[224]), .outData_225(wire_switch_out_stage6[225]), .outData_226(wire_switch_out_stage6[226]), .outData_227(wire_switch_out_stage6[227]), .outData_228(wire_switch_out_stage6[228]), .outData_229(wire_switch_out_stage6[229]), .outData_230(wire_switch_out_stage6[230]), .outData_231(wire_switch_out_stage6[231]), .outData_232(wire_switch_out_stage6[232]), .outData_233(wire_switch_out_stage6[233]), .outData_234(wire_switch_out_stage6[234]), .outData_235(wire_switch_out_stage6[235]), .outData_236(wire_switch_out_stage6[236]), .outData_237(wire_switch_out_stage6[237]), .outData_238(wire_switch_out_stage6[238]), .outData_239(wire_switch_out_stage6[239]), .outData_240(wire_switch_out_stage6[240]), .outData_241(wire_switch_out_stage6[241]), .outData_242(wire_switch_out_stage6[242]), .outData_243(wire_switch_out_stage6[243]), .outData_244(wire_switch_out_stage6[244]), .outData_245(wire_switch_out_stage6[245]), .outData_246(wire_switch_out_stage6[246]), .outData_247(wire_switch_out_stage6[247]), .outData_248(wire_switch_out_stage6[248]), .outData_249(wire_switch_out_stage6[249]), .outData_250(wire_switch_out_stage6[250]), .outData_251(wire_switch_out_stage6[251]), .outData_252(wire_switch_out_stage6[252]), .outData_253(wire_switch_out_stage6[253]), .outData_254(wire_switch_out_stage6[254]), .outData_255(wire_switch_out_stage6[255]), 
        .in_start(con_in_start_stage6), .out_start(in_start_stage5), .ctrl(wire_ctrl_stage6), .clk(clk), .rst(rst));
  
  wireCon_dp256_st6_R wire_stage_6(
        .inData_0(wire_switch_out_stage7[0]), .inData_1(wire_switch_out_stage7[1]), .inData_2(wire_switch_out_stage7[2]), .inData_3(wire_switch_out_stage7[3]), .inData_4(wire_switch_out_stage7[4]), .inData_5(wire_switch_out_stage7[5]), .inData_6(wire_switch_out_stage7[6]), .inData_7(wire_switch_out_stage7[7]), .inData_8(wire_switch_out_stage7[8]), .inData_9(wire_switch_out_stage7[9]), .inData_10(wire_switch_out_stage7[10]), .inData_11(wire_switch_out_stage7[11]), .inData_12(wire_switch_out_stage7[12]), .inData_13(wire_switch_out_stage7[13]), .inData_14(wire_switch_out_stage7[14]), .inData_15(wire_switch_out_stage7[15]), .inData_16(wire_switch_out_stage7[16]), .inData_17(wire_switch_out_stage7[17]), .inData_18(wire_switch_out_stage7[18]), .inData_19(wire_switch_out_stage7[19]), .inData_20(wire_switch_out_stage7[20]), .inData_21(wire_switch_out_stage7[21]), .inData_22(wire_switch_out_stage7[22]), .inData_23(wire_switch_out_stage7[23]), .inData_24(wire_switch_out_stage7[24]), .inData_25(wire_switch_out_stage7[25]), .inData_26(wire_switch_out_stage7[26]), .inData_27(wire_switch_out_stage7[27]), .inData_28(wire_switch_out_stage7[28]), .inData_29(wire_switch_out_stage7[29]), .inData_30(wire_switch_out_stage7[30]), .inData_31(wire_switch_out_stage7[31]), .inData_32(wire_switch_out_stage7[32]), .inData_33(wire_switch_out_stage7[33]), .inData_34(wire_switch_out_stage7[34]), .inData_35(wire_switch_out_stage7[35]), .inData_36(wire_switch_out_stage7[36]), .inData_37(wire_switch_out_stage7[37]), .inData_38(wire_switch_out_stage7[38]), .inData_39(wire_switch_out_stage7[39]), .inData_40(wire_switch_out_stage7[40]), .inData_41(wire_switch_out_stage7[41]), .inData_42(wire_switch_out_stage7[42]), .inData_43(wire_switch_out_stage7[43]), .inData_44(wire_switch_out_stage7[44]), .inData_45(wire_switch_out_stage7[45]), .inData_46(wire_switch_out_stage7[46]), .inData_47(wire_switch_out_stage7[47]), .inData_48(wire_switch_out_stage7[48]), .inData_49(wire_switch_out_stage7[49]), .inData_50(wire_switch_out_stage7[50]), .inData_51(wire_switch_out_stage7[51]), .inData_52(wire_switch_out_stage7[52]), .inData_53(wire_switch_out_stage7[53]), .inData_54(wire_switch_out_stage7[54]), .inData_55(wire_switch_out_stage7[55]), .inData_56(wire_switch_out_stage7[56]), .inData_57(wire_switch_out_stage7[57]), .inData_58(wire_switch_out_stage7[58]), .inData_59(wire_switch_out_stage7[59]), .inData_60(wire_switch_out_stage7[60]), .inData_61(wire_switch_out_stage7[61]), .inData_62(wire_switch_out_stage7[62]), .inData_63(wire_switch_out_stage7[63]), .inData_64(wire_switch_out_stage7[64]), .inData_65(wire_switch_out_stage7[65]), .inData_66(wire_switch_out_stage7[66]), .inData_67(wire_switch_out_stage7[67]), .inData_68(wire_switch_out_stage7[68]), .inData_69(wire_switch_out_stage7[69]), .inData_70(wire_switch_out_stage7[70]), .inData_71(wire_switch_out_stage7[71]), .inData_72(wire_switch_out_stage7[72]), .inData_73(wire_switch_out_stage7[73]), .inData_74(wire_switch_out_stage7[74]), .inData_75(wire_switch_out_stage7[75]), .inData_76(wire_switch_out_stage7[76]), .inData_77(wire_switch_out_stage7[77]), .inData_78(wire_switch_out_stage7[78]), .inData_79(wire_switch_out_stage7[79]), .inData_80(wire_switch_out_stage7[80]), .inData_81(wire_switch_out_stage7[81]), .inData_82(wire_switch_out_stage7[82]), .inData_83(wire_switch_out_stage7[83]), .inData_84(wire_switch_out_stage7[84]), .inData_85(wire_switch_out_stage7[85]), .inData_86(wire_switch_out_stage7[86]), .inData_87(wire_switch_out_stage7[87]), .inData_88(wire_switch_out_stage7[88]), .inData_89(wire_switch_out_stage7[89]), .inData_90(wire_switch_out_stage7[90]), .inData_91(wire_switch_out_stage7[91]), .inData_92(wire_switch_out_stage7[92]), .inData_93(wire_switch_out_stage7[93]), .inData_94(wire_switch_out_stage7[94]), .inData_95(wire_switch_out_stage7[95]), .inData_96(wire_switch_out_stage7[96]), .inData_97(wire_switch_out_stage7[97]), .inData_98(wire_switch_out_stage7[98]), .inData_99(wire_switch_out_stage7[99]), .inData_100(wire_switch_out_stage7[100]), .inData_101(wire_switch_out_stage7[101]), .inData_102(wire_switch_out_stage7[102]), .inData_103(wire_switch_out_stage7[103]), .inData_104(wire_switch_out_stage7[104]), .inData_105(wire_switch_out_stage7[105]), .inData_106(wire_switch_out_stage7[106]), .inData_107(wire_switch_out_stage7[107]), .inData_108(wire_switch_out_stage7[108]), .inData_109(wire_switch_out_stage7[109]), .inData_110(wire_switch_out_stage7[110]), .inData_111(wire_switch_out_stage7[111]), .inData_112(wire_switch_out_stage7[112]), .inData_113(wire_switch_out_stage7[113]), .inData_114(wire_switch_out_stage7[114]), .inData_115(wire_switch_out_stage7[115]), .inData_116(wire_switch_out_stage7[116]), .inData_117(wire_switch_out_stage7[117]), .inData_118(wire_switch_out_stage7[118]), .inData_119(wire_switch_out_stage7[119]), .inData_120(wire_switch_out_stage7[120]), .inData_121(wire_switch_out_stage7[121]), .inData_122(wire_switch_out_stage7[122]), .inData_123(wire_switch_out_stage7[123]), .inData_124(wire_switch_out_stage7[124]), .inData_125(wire_switch_out_stage7[125]), .inData_126(wire_switch_out_stage7[126]), .inData_127(wire_switch_out_stage7[127]), .inData_128(wire_switch_out_stage7[128]), .inData_129(wire_switch_out_stage7[129]), .inData_130(wire_switch_out_stage7[130]), .inData_131(wire_switch_out_stage7[131]), .inData_132(wire_switch_out_stage7[132]), .inData_133(wire_switch_out_stage7[133]), .inData_134(wire_switch_out_stage7[134]), .inData_135(wire_switch_out_stage7[135]), .inData_136(wire_switch_out_stage7[136]), .inData_137(wire_switch_out_stage7[137]), .inData_138(wire_switch_out_stage7[138]), .inData_139(wire_switch_out_stage7[139]), .inData_140(wire_switch_out_stage7[140]), .inData_141(wire_switch_out_stage7[141]), .inData_142(wire_switch_out_stage7[142]), .inData_143(wire_switch_out_stage7[143]), .inData_144(wire_switch_out_stage7[144]), .inData_145(wire_switch_out_stage7[145]), .inData_146(wire_switch_out_stage7[146]), .inData_147(wire_switch_out_stage7[147]), .inData_148(wire_switch_out_stage7[148]), .inData_149(wire_switch_out_stage7[149]), .inData_150(wire_switch_out_stage7[150]), .inData_151(wire_switch_out_stage7[151]), .inData_152(wire_switch_out_stage7[152]), .inData_153(wire_switch_out_stage7[153]), .inData_154(wire_switch_out_stage7[154]), .inData_155(wire_switch_out_stage7[155]), .inData_156(wire_switch_out_stage7[156]), .inData_157(wire_switch_out_stage7[157]), .inData_158(wire_switch_out_stage7[158]), .inData_159(wire_switch_out_stage7[159]), .inData_160(wire_switch_out_stage7[160]), .inData_161(wire_switch_out_stage7[161]), .inData_162(wire_switch_out_stage7[162]), .inData_163(wire_switch_out_stage7[163]), .inData_164(wire_switch_out_stage7[164]), .inData_165(wire_switch_out_stage7[165]), .inData_166(wire_switch_out_stage7[166]), .inData_167(wire_switch_out_stage7[167]), .inData_168(wire_switch_out_stage7[168]), .inData_169(wire_switch_out_stage7[169]), .inData_170(wire_switch_out_stage7[170]), .inData_171(wire_switch_out_stage7[171]), .inData_172(wire_switch_out_stage7[172]), .inData_173(wire_switch_out_stage7[173]), .inData_174(wire_switch_out_stage7[174]), .inData_175(wire_switch_out_stage7[175]), .inData_176(wire_switch_out_stage7[176]), .inData_177(wire_switch_out_stage7[177]), .inData_178(wire_switch_out_stage7[178]), .inData_179(wire_switch_out_stage7[179]), .inData_180(wire_switch_out_stage7[180]), .inData_181(wire_switch_out_stage7[181]), .inData_182(wire_switch_out_stage7[182]), .inData_183(wire_switch_out_stage7[183]), .inData_184(wire_switch_out_stage7[184]), .inData_185(wire_switch_out_stage7[185]), .inData_186(wire_switch_out_stage7[186]), .inData_187(wire_switch_out_stage7[187]), .inData_188(wire_switch_out_stage7[188]), .inData_189(wire_switch_out_stage7[189]), .inData_190(wire_switch_out_stage7[190]), .inData_191(wire_switch_out_stage7[191]), .inData_192(wire_switch_out_stage7[192]), .inData_193(wire_switch_out_stage7[193]), .inData_194(wire_switch_out_stage7[194]), .inData_195(wire_switch_out_stage7[195]), .inData_196(wire_switch_out_stage7[196]), .inData_197(wire_switch_out_stage7[197]), .inData_198(wire_switch_out_stage7[198]), .inData_199(wire_switch_out_stage7[199]), .inData_200(wire_switch_out_stage7[200]), .inData_201(wire_switch_out_stage7[201]), .inData_202(wire_switch_out_stage7[202]), .inData_203(wire_switch_out_stage7[203]), .inData_204(wire_switch_out_stage7[204]), .inData_205(wire_switch_out_stage7[205]), .inData_206(wire_switch_out_stage7[206]), .inData_207(wire_switch_out_stage7[207]), .inData_208(wire_switch_out_stage7[208]), .inData_209(wire_switch_out_stage7[209]), .inData_210(wire_switch_out_stage7[210]), .inData_211(wire_switch_out_stage7[211]), .inData_212(wire_switch_out_stage7[212]), .inData_213(wire_switch_out_stage7[213]), .inData_214(wire_switch_out_stage7[214]), .inData_215(wire_switch_out_stage7[215]), .inData_216(wire_switch_out_stage7[216]), .inData_217(wire_switch_out_stage7[217]), .inData_218(wire_switch_out_stage7[218]), .inData_219(wire_switch_out_stage7[219]), .inData_220(wire_switch_out_stage7[220]), .inData_221(wire_switch_out_stage7[221]), .inData_222(wire_switch_out_stage7[222]), .inData_223(wire_switch_out_stage7[223]), .inData_224(wire_switch_out_stage7[224]), .inData_225(wire_switch_out_stage7[225]), .inData_226(wire_switch_out_stage7[226]), .inData_227(wire_switch_out_stage7[227]), .inData_228(wire_switch_out_stage7[228]), .inData_229(wire_switch_out_stage7[229]), .inData_230(wire_switch_out_stage7[230]), .inData_231(wire_switch_out_stage7[231]), .inData_232(wire_switch_out_stage7[232]), .inData_233(wire_switch_out_stage7[233]), .inData_234(wire_switch_out_stage7[234]), .inData_235(wire_switch_out_stage7[235]), .inData_236(wire_switch_out_stage7[236]), .inData_237(wire_switch_out_stage7[237]), .inData_238(wire_switch_out_stage7[238]), .inData_239(wire_switch_out_stage7[239]), .inData_240(wire_switch_out_stage7[240]), .inData_241(wire_switch_out_stage7[241]), .inData_242(wire_switch_out_stage7[242]), .inData_243(wire_switch_out_stage7[243]), .inData_244(wire_switch_out_stage7[244]), .inData_245(wire_switch_out_stage7[245]), .inData_246(wire_switch_out_stage7[246]), .inData_247(wire_switch_out_stage7[247]), .inData_248(wire_switch_out_stage7[248]), .inData_249(wire_switch_out_stage7[249]), .inData_250(wire_switch_out_stage7[250]), .inData_251(wire_switch_out_stage7[251]), .inData_252(wire_switch_out_stage7[252]), .inData_253(wire_switch_out_stage7[253]), .inData_254(wire_switch_out_stage7[254]), .inData_255(wire_switch_out_stage7[255]), 
        .outData_0(wire_switch_in_stage6[0]), .outData_1(wire_switch_in_stage6[1]), .outData_2(wire_switch_in_stage6[2]), .outData_3(wire_switch_in_stage6[3]), .outData_4(wire_switch_in_stage6[4]), .outData_5(wire_switch_in_stage6[5]), .outData_6(wire_switch_in_stage6[6]), .outData_7(wire_switch_in_stage6[7]), .outData_8(wire_switch_in_stage6[8]), .outData_9(wire_switch_in_stage6[9]), .outData_10(wire_switch_in_stage6[10]), .outData_11(wire_switch_in_stage6[11]), .outData_12(wire_switch_in_stage6[12]), .outData_13(wire_switch_in_stage6[13]), .outData_14(wire_switch_in_stage6[14]), .outData_15(wire_switch_in_stage6[15]), .outData_16(wire_switch_in_stage6[16]), .outData_17(wire_switch_in_stage6[17]), .outData_18(wire_switch_in_stage6[18]), .outData_19(wire_switch_in_stage6[19]), .outData_20(wire_switch_in_stage6[20]), .outData_21(wire_switch_in_stage6[21]), .outData_22(wire_switch_in_stage6[22]), .outData_23(wire_switch_in_stage6[23]), .outData_24(wire_switch_in_stage6[24]), .outData_25(wire_switch_in_stage6[25]), .outData_26(wire_switch_in_stage6[26]), .outData_27(wire_switch_in_stage6[27]), .outData_28(wire_switch_in_stage6[28]), .outData_29(wire_switch_in_stage6[29]), .outData_30(wire_switch_in_stage6[30]), .outData_31(wire_switch_in_stage6[31]), .outData_32(wire_switch_in_stage6[32]), .outData_33(wire_switch_in_stage6[33]), .outData_34(wire_switch_in_stage6[34]), .outData_35(wire_switch_in_stage6[35]), .outData_36(wire_switch_in_stage6[36]), .outData_37(wire_switch_in_stage6[37]), .outData_38(wire_switch_in_stage6[38]), .outData_39(wire_switch_in_stage6[39]), .outData_40(wire_switch_in_stage6[40]), .outData_41(wire_switch_in_stage6[41]), .outData_42(wire_switch_in_stage6[42]), .outData_43(wire_switch_in_stage6[43]), .outData_44(wire_switch_in_stage6[44]), .outData_45(wire_switch_in_stage6[45]), .outData_46(wire_switch_in_stage6[46]), .outData_47(wire_switch_in_stage6[47]), .outData_48(wire_switch_in_stage6[48]), .outData_49(wire_switch_in_stage6[49]), .outData_50(wire_switch_in_stage6[50]), .outData_51(wire_switch_in_stage6[51]), .outData_52(wire_switch_in_stage6[52]), .outData_53(wire_switch_in_stage6[53]), .outData_54(wire_switch_in_stage6[54]), .outData_55(wire_switch_in_stage6[55]), .outData_56(wire_switch_in_stage6[56]), .outData_57(wire_switch_in_stage6[57]), .outData_58(wire_switch_in_stage6[58]), .outData_59(wire_switch_in_stage6[59]), .outData_60(wire_switch_in_stage6[60]), .outData_61(wire_switch_in_stage6[61]), .outData_62(wire_switch_in_stage6[62]), .outData_63(wire_switch_in_stage6[63]), .outData_64(wire_switch_in_stage6[64]), .outData_65(wire_switch_in_stage6[65]), .outData_66(wire_switch_in_stage6[66]), .outData_67(wire_switch_in_stage6[67]), .outData_68(wire_switch_in_stage6[68]), .outData_69(wire_switch_in_stage6[69]), .outData_70(wire_switch_in_stage6[70]), .outData_71(wire_switch_in_stage6[71]), .outData_72(wire_switch_in_stage6[72]), .outData_73(wire_switch_in_stage6[73]), .outData_74(wire_switch_in_stage6[74]), .outData_75(wire_switch_in_stage6[75]), .outData_76(wire_switch_in_stage6[76]), .outData_77(wire_switch_in_stage6[77]), .outData_78(wire_switch_in_stage6[78]), .outData_79(wire_switch_in_stage6[79]), .outData_80(wire_switch_in_stage6[80]), .outData_81(wire_switch_in_stage6[81]), .outData_82(wire_switch_in_stage6[82]), .outData_83(wire_switch_in_stage6[83]), .outData_84(wire_switch_in_stage6[84]), .outData_85(wire_switch_in_stage6[85]), .outData_86(wire_switch_in_stage6[86]), .outData_87(wire_switch_in_stage6[87]), .outData_88(wire_switch_in_stage6[88]), .outData_89(wire_switch_in_stage6[89]), .outData_90(wire_switch_in_stage6[90]), .outData_91(wire_switch_in_stage6[91]), .outData_92(wire_switch_in_stage6[92]), .outData_93(wire_switch_in_stage6[93]), .outData_94(wire_switch_in_stage6[94]), .outData_95(wire_switch_in_stage6[95]), .outData_96(wire_switch_in_stage6[96]), .outData_97(wire_switch_in_stage6[97]), .outData_98(wire_switch_in_stage6[98]), .outData_99(wire_switch_in_stage6[99]), .outData_100(wire_switch_in_stage6[100]), .outData_101(wire_switch_in_stage6[101]), .outData_102(wire_switch_in_stage6[102]), .outData_103(wire_switch_in_stage6[103]), .outData_104(wire_switch_in_stage6[104]), .outData_105(wire_switch_in_stage6[105]), .outData_106(wire_switch_in_stage6[106]), .outData_107(wire_switch_in_stage6[107]), .outData_108(wire_switch_in_stage6[108]), .outData_109(wire_switch_in_stage6[109]), .outData_110(wire_switch_in_stage6[110]), .outData_111(wire_switch_in_stage6[111]), .outData_112(wire_switch_in_stage6[112]), .outData_113(wire_switch_in_stage6[113]), .outData_114(wire_switch_in_stage6[114]), .outData_115(wire_switch_in_stage6[115]), .outData_116(wire_switch_in_stage6[116]), .outData_117(wire_switch_in_stage6[117]), .outData_118(wire_switch_in_stage6[118]), .outData_119(wire_switch_in_stage6[119]), .outData_120(wire_switch_in_stage6[120]), .outData_121(wire_switch_in_stage6[121]), .outData_122(wire_switch_in_stage6[122]), .outData_123(wire_switch_in_stage6[123]), .outData_124(wire_switch_in_stage6[124]), .outData_125(wire_switch_in_stage6[125]), .outData_126(wire_switch_in_stage6[126]), .outData_127(wire_switch_in_stage6[127]), .outData_128(wire_switch_in_stage6[128]), .outData_129(wire_switch_in_stage6[129]), .outData_130(wire_switch_in_stage6[130]), .outData_131(wire_switch_in_stage6[131]), .outData_132(wire_switch_in_stage6[132]), .outData_133(wire_switch_in_stage6[133]), .outData_134(wire_switch_in_stage6[134]), .outData_135(wire_switch_in_stage6[135]), .outData_136(wire_switch_in_stage6[136]), .outData_137(wire_switch_in_stage6[137]), .outData_138(wire_switch_in_stage6[138]), .outData_139(wire_switch_in_stage6[139]), .outData_140(wire_switch_in_stage6[140]), .outData_141(wire_switch_in_stage6[141]), .outData_142(wire_switch_in_stage6[142]), .outData_143(wire_switch_in_stage6[143]), .outData_144(wire_switch_in_stage6[144]), .outData_145(wire_switch_in_stage6[145]), .outData_146(wire_switch_in_stage6[146]), .outData_147(wire_switch_in_stage6[147]), .outData_148(wire_switch_in_stage6[148]), .outData_149(wire_switch_in_stage6[149]), .outData_150(wire_switch_in_stage6[150]), .outData_151(wire_switch_in_stage6[151]), .outData_152(wire_switch_in_stage6[152]), .outData_153(wire_switch_in_stage6[153]), .outData_154(wire_switch_in_stage6[154]), .outData_155(wire_switch_in_stage6[155]), .outData_156(wire_switch_in_stage6[156]), .outData_157(wire_switch_in_stage6[157]), .outData_158(wire_switch_in_stage6[158]), .outData_159(wire_switch_in_stage6[159]), .outData_160(wire_switch_in_stage6[160]), .outData_161(wire_switch_in_stage6[161]), .outData_162(wire_switch_in_stage6[162]), .outData_163(wire_switch_in_stage6[163]), .outData_164(wire_switch_in_stage6[164]), .outData_165(wire_switch_in_stage6[165]), .outData_166(wire_switch_in_stage6[166]), .outData_167(wire_switch_in_stage6[167]), .outData_168(wire_switch_in_stage6[168]), .outData_169(wire_switch_in_stage6[169]), .outData_170(wire_switch_in_stage6[170]), .outData_171(wire_switch_in_stage6[171]), .outData_172(wire_switch_in_stage6[172]), .outData_173(wire_switch_in_stage6[173]), .outData_174(wire_switch_in_stage6[174]), .outData_175(wire_switch_in_stage6[175]), .outData_176(wire_switch_in_stage6[176]), .outData_177(wire_switch_in_stage6[177]), .outData_178(wire_switch_in_stage6[178]), .outData_179(wire_switch_in_stage6[179]), .outData_180(wire_switch_in_stage6[180]), .outData_181(wire_switch_in_stage6[181]), .outData_182(wire_switch_in_stage6[182]), .outData_183(wire_switch_in_stage6[183]), .outData_184(wire_switch_in_stage6[184]), .outData_185(wire_switch_in_stage6[185]), .outData_186(wire_switch_in_stage6[186]), .outData_187(wire_switch_in_stage6[187]), .outData_188(wire_switch_in_stage6[188]), .outData_189(wire_switch_in_stage6[189]), .outData_190(wire_switch_in_stage6[190]), .outData_191(wire_switch_in_stage6[191]), .outData_192(wire_switch_in_stage6[192]), .outData_193(wire_switch_in_stage6[193]), .outData_194(wire_switch_in_stage6[194]), .outData_195(wire_switch_in_stage6[195]), .outData_196(wire_switch_in_stage6[196]), .outData_197(wire_switch_in_stage6[197]), .outData_198(wire_switch_in_stage6[198]), .outData_199(wire_switch_in_stage6[199]), .outData_200(wire_switch_in_stage6[200]), .outData_201(wire_switch_in_stage6[201]), .outData_202(wire_switch_in_stage6[202]), .outData_203(wire_switch_in_stage6[203]), .outData_204(wire_switch_in_stage6[204]), .outData_205(wire_switch_in_stage6[205]), .outData_206(wire_switch_in_stage6[206]), .outData_207(wire_switch_in_stage6[207]), .outData_208(wire_switch_in_stage6[208]), .outData_209(wire_switch_in_stage6[209]), .outData_210(wire_switch_in_stage6[210]), .outData_211(wire_switch_in_stage6[211]), .outData_212(wire_switch_in_stage6[212]), .outData_213(wire_switch_in_stage6[213]), .outData_214(wire_switch_in_stage6[214]), .outData_215(wire_switch_in_stage6[215]), .outData_216(wire_switch_in_stage6[216]), .outData_217(wire_switch_in_stage6[217]), .outData_218(wire_switch_in_stage6[218]), .outData_219(wire_switch_in_stage6[219]), .outData_220(wire_switch_in_stage6[220]), .outData_221(wire_switch_in_stage6[221]), .outData_222(wire_switch_in_stage6[222]), .outData_223(wire_switch_in_stage6[223]), .outData_224(wire_switch_in_stage6[224]), .outData_225(wire_switch_in_stage6[225]), .outData_226(wire_switch_in_stage6[226]), .outData_227(wire_switch_in_stage6[227]), .outData_228(wire_switch_in_stage6[228]), .outData_229(wire_switch_in_stage6[229]), .outData_230(wire_switch_in_stage6[230]), .outData_231(wire_switch_in_stage6[231]), .outData_232(wire_switch_in_stage6[232]), .outData_233(wire_switch_in_stage6[233]), .outData_234(wire_switch_in_stage6[234]), .outData_235(wire_switch_in_stage6[235]), .outData_236(wire_switch_in_stage6[236]), .outData_237(wire_switch_in_stage6[237]), .outData_238(wire_switch_in_stage6[238]), .outData_239(wire_switch_in_stage6[239]), .outData_240(wire_switch_in_stage6[240]), .outData_241(wire_switch_in_stage6[241]), .outData_242(wire_switch_in_stage6[242]), .outData_243(wire_switch_in_stage6[243]), .outData_244(wire_switch_in_stage6[244]), .outData_245(wire_switch_in_stage6[245]), .outData_246(wire_switch_in_stage6[246]), .outData_247(wire_switch_in_stage6[247]), .outData_248(wire_switch_in_stage6[248]), .outData_249(wire_switch_in_stage6[249]), .outData_250(wire_switch_in_stage6[250]), .outData_251(wire_switch_in_stage6[251]), .outData_252(wire_switch_in_stage6[252]), .outData_253(wire_switch_in_stage6[253]), .outData_254(wire_switch_in_stage6[254]), .outData_255(wire_switch_in_stage6[255]), 
        .in_start(in_start_stage6), .out_start(con_in_start_stage6), .clk(clk), .rst(rst)); 

  
  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[0] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[1] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[2] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[3] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[4] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[5] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[6] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[7] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[8] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[9] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[10] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[11] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[12] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[13] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[14] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[15] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[16] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[17] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[18] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[19] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[20] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[21] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[22] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[23] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[24] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[25] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[26] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[27] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[28] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[29] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[30] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[31] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[32] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[33] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[34] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[35] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[36] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[37] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[38] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[39] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[40] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[41] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[42] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[43] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[44] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[45] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[46] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[47] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[48] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[49] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[50] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[51] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[52] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[53] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[54] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[55] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[56] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[57] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[58] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[59] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[60] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[61] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[62] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[63] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[64] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[65] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[66] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[67] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[68] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[69] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[70] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[71] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[72] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[73] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[74] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[75] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[76] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[77] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[78] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[79] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[80] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[81] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[82] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[83] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[84] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[85] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[86] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[87] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[88] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[89] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[90] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[91] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[92] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[93] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[94] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[95] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[96] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[97] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[98] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[99] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[100] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[101] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[102] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[103] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[104] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[105] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[106] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[107] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[108] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[109] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[110] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[111] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[112] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[113] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[114] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[115] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[116] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[117] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[118] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[119] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[120] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[121] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[122] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[123] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[124] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[125] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[126] <= counter_w[1]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage6[127] <= counter_w[1]; 
  end                            

  wire [DATA_WIDTH-1:0] wire_switch_in_stage5[255:0];
  wire [DATA_WIDTH-1:0] wire_switch_out_stage5[255:0];
  reg [127:0] wire_ctrl_stage5;

  switches_stage_st5_0_R switch_stage_5(
        .inData_0(wire_switch_in_stage5[0]), .inData_1(wire_switch_in_stage5[1]), .inData_2(wire_switch_in_stage5[2]), .inData_3(wire_switch_in_stage5[3]), .inData_4(wire_switch_in_stage5[4]), .inData_5(wire_switch_in_stage5[5]), .inData_6(wire_switch_in_stage5[6]), .inData_7(wire_switch_in_stage5[7]), .inData_8(wire_switch_in_stage5[8]), .inData_9(wire_switch_in_stage5[9]), .inData_10(wire_switch_in_stage5[10]), .inData_11(wire_switch_in_stage5[11]), .inData_12(wire_switch_in_stage5[12]), .inData_13(wire_switch_in_stage5[13]), .inData_14(wire_switch_in_stage5[14]), .inData_15(wire_switch_in_stage5[15]), .inData_16(wire_switch_in_stage5[16]), .inData_17(wire_switch_in_stage5[17]), .inData_18(wire_switch_in_stage5[18]), .inData_19(wire_switch_in_stage5[19]), .inData_20(wire_switch_in_stage5[20]), .inData_21(wire_switch_in_stage5[21]), .inData_22(wire_switch_in_stage5[22]), .inData_23(wire_switch_in_stage5[23]), .inData_24(wire_switch_in_stage5[24]), .inData_25(wire_switch_in_stage5[25]), .inData_26(wire_switch_in_stage5[26]), .inData_27(wire_switch_in_stage5[27]), .inData_28(wire_switch_in_stage5[28]), .inData_29(wire_switch_in_stage5[29]), .inData_30(wire_switch_in_stage5[30]), .inData_31(wire_switch_in_stage5[31]), .inData_32(wire_switch_in_stage5[32]), .inData_33(wire_switch_in_stage5[33]), .inData_34(wire_switch_in_stage5[34]), .inData_35(wire_switch_in_stage5[35]), .inData_36(wire_switch_in_stage5[36]), .inData_37(wire_switch_in_stage5[37]), .inData_38(wire_switch_in_stage5[38]), .inData_39(wire_switch_in_stage5[39]), .inData_40(wire_switch_in_stage5[40]), .inData_41(wire_switch_in_stage5[41]), .inData_42(wire_switch_in_stage5[42]), .inData_43(wire_switch_in_stage5[43]), .inData_44(wire_switch_in_stage5[44]), .inData_45(wire_switch_in_stage5[45]), .inData_46(wire_switch_in_stage5[46]), .inData_47(wire_switch_in_stage5[47]), .inData_48(wire_switch_in_stage5[48]), .inData_49(wire_switch_in_stage5[49]), .inData_50(wire_switch_in_stage5[50]), .inData_51(wire_switch_in_stage5[51]), .inData_52(wire_switch_in_stage5[52]), .inData_53(wire_switch_in_stage5[53]), .inData_54(wire_switch_in_stage5[54]), .inData_55(wire_switch_in_stage5[55]), .inData_56(wire_switch_in_stage5[56]), .inData_57(wire_switch_in_stage5[57]), .inData_58(wire_switch_in_stage5[58]), .inData_59(wire_switch_in_stage5[59]), .inData_60(wire_switch_in_stage5[60]), .inData_61(wire_switch_in_stage5[61]), .inData_62(wire_switch_in_stage5[62]), .inData_63(wire_switch_in_stage5[63]), .inData_64(wire_switch_in_stage5[64]), .inData_65(wire_switch_in_stage5[65]), .inData_66(wire_switch_in_stage5[66]), .inData_67(wire_switch_in_stage5[67]), .inData_68(wire_switch_in_stage5[68]), .inData_69(wire_switch_in_stage5[69]), .inData_70(wire_switch_in_stage5[70]), .inData_71(wire_switch_in_stage5[71]), .inData_72(wire_switch_in_stage5[72]), .inData_73(wire_switch_in_stage5[73]), .inData_74(wire_switch_in_stage5[74]), .inData_75(wire_switch_in_stage5[75]), .inData_76(wire_switch_in_stage5[76]), .inData_77(wire_switch_in_stage5[77]), .inData_78(wire_switch_in_stage5[78]), .inData_79(wire_switch_in_stage5[79]), .inData_80(wire_switch_in_stage5[80]), .inData_81(wire_switch_in_stage5[81]), .inData_82(wire_switch_in_stage5[82]), .inData_83(wire_switch_in_stage5[83]), .inData_84(wire_switch_in_stage5[84]), .inData_85(wire_switch_in_stage5[85]), .inData_86(wire_switch_in_stage5[86]), .inData_87(wire_switch_in_stage5[87]), .inData_88(wire_switch_in_stage5[88]), .inData_89(wire_switch_in_stage5[89]), .inData_90(wire_switch_in_stage5[90]), .inData_91(wire_switch_in_stage5[91]), .inData_92(wire_switch_in_stage5[92]), .inData_93(wire_switch_in_stage5[93]), .inData_94(wire_switch_in_stage5[94]), .inData_95(wire_switch_in_stage5[95]), .inData_96(wire_switch_in_stage5[96]), .inData_97(wire_switch_in_stage5[97]), .inData_98(wire_switch_in_stage5[98]), .inData_99(wire_switch_in_stage5[99]), .inData_100(wire_switch_in_stage5[100]), .inData_101(wire_switch_in_stage5[101]), .inData_102(wire_switch_in_stage5[102]), .inData_103(wire_switch_in_stage5[103]), .inData_104(wire_switch_in_stage5[104]), .inData_105(wire_switch_in_stage5[105]), .inData_106(wire_switch_in_stage5[106]), .inData_107(wire_switch_in_stage5[107]), .inData_108(wire_switch_in_stage5[108]), .inData_109(wire_switch_in_stage5[109]), .inData_110(wire_switch_in_stage5[110]), .inData_111(wire_switch_in_stage5[111]), .inData_112(wire_switch_in_stage5[112]), .inData_113(wire_switch_in_stage5[113]), .inData_114(wire_switch_in_stage5[114]), .inData_115(wire_switch_in_stage5[115]), .inData_116(wire_switch_in_stage5[116]), .inData_117(wire_switch_in_stage5[117]), .inData_118(wire_switch_in_stage5[118]), .inData_119(wire_switch_in_stage5[119]), .inData_120(wire_switch_in_stage5[120]), .inData_121(wire_switch_in_stage5[121]), .inData_122(wire_switch_in_stage5[122]), .inData_123(wire_switch_in_stage5[123]), .inData_124(wire_switch_in_stage5[124]), .inData_125(wire_switch_in_stage5[125]), .inData_126(wire_switch_in_stage5[126]), .inData_127(wire_switch_in_stage5[127]), .inData_128(wire_switch_in_stage5[128]), .inData_129(wire_switch_in_stage5[129]), .inData_130(wire_switch_in_stage5[130]), .inData_131(wire_switch_in_stage5[131]), .inData_132(wire_switch_in_stage5[132]), .inData_133(wire_switch_in_stage5[133]), .inData_134(wire_switch_in_stage5[134]), .inData_135(wire_switch_in_stage5[135]), .inData_136(wire_switch_in_stage5[136]), .inData_137(wire_switch_in_stage5[137]), .inData_138(wire_switch_in_stage5[138]), .inData_139(wire_switch_in_stage5[139]), .inData_140(wire_switch_in_stage5[140]), .inData_141(wire_switch_in_stage5[141]), .inData_142(wire_switch_in_stage5[142]), .inData_143(wire_switch_in_stage5[143]), .inData_144(wire_switch_in_stage5[144]), .inData_145(wire_switch_in_stage5[145]), .inData_146(wire_switch_in_stage5[146]), .inData_147(wire_switch_in_stage5[147]), .inData_148(wire_switch_in_stage5[148]), .inData_149(wire_switch_in_stage5[149]), .inData_150(wire_switch_in_stage5[150]), .inData_151(wire_switch_in_stage5[151]), .inData_152(wire_switch_in_stage5[152]), .inData_153(wire_switch_in_stage5[153]), .inData_154(wire_switch_in_stage5[154]), .inData_155(wire_switch_in_stage5[155]), .inData_156(wire_switch_in_stage5[156]), .inData_157(wire_switch_in_stage5[157]), .inData_158(wire_switch_in_stage5[158]), .inData_159(wire_switch_in_stage5[159]), .inData_160(wire_switch_in_stage5[160]), .inData_161(wire_switch_in_stage5[161]), .inData_162(wire_switch_in_stage5[162]), .inData_163(wire_switch_in_stage5[163]), .inData_164(wire_switch_in_stage5[164]), .inData_165(wire_switch_in_stage5[165]), .inData_166(wire_switch_in_stage5[166]), .inData_167(wire_switch_in_stage5[167]), .inData_168(wire_switch_in_stage5[168]), .inData_169(wire_switch_in_stage5[169]), .inData_170(wire_switch_in_stage5[170]), .inData_171(wire_switch_in_stage5[171]), .inData_172(wire_switch_in_stage5[172]), .inData_173(wire_switch_in_stage5[173]), .inData_174(wire_switch_in_stage5[174]), .inData_175(wire_switch_in_stage5[175]), .inData_176(wire_switch_in_stage5[176]), .inData_177(wire_switch_in_stage5[177]), .inData_178(wire_switch_in_stage5[178]), .inData_179(wire_switch_in_stage5[179]), .inData_180(wire_switch_in_stage5[180]), .inData_181(wire_switch_in_stage5[181]), .inData_182(wire_switch_in_stage5[182]), .inData_183(wire_switch_in_stage5[183]), .inData_184(wire_switch_in_stage5[184]), .inData_185(wire_switch_in_stage5[185]), .inData_186(wire_switch_in_stage5[186]), .inData_187(wire_switch_in_stage5[187]), .inData_188(wire_switch_in_stage5[188]), .inData_189(wire_switch_in_stage5[189]), .inData_190(wire_switch_in_stage5[190]), .inData_191(wire_switch_in_stage5[191]), .inData_192(wire_switch_in_stage5[192]), .inData_193(wire_switch_in_stage5[193]), .inData_194(wire_switch_in_stage5[194]), .inData_195(wire_switch_in_stage5[195]), .inData_196(wire_switch_in_stage5[196]), .inData_197(wire_switch_in_stage5[197]), .inData_198(wire_switch_in_stage5[198]), .inData_199(wire_switch_in_stage5[199]), .inData_200(wire_switch_in_stage5[200]), .inData_201(wire_switch_in_stage5[201]), .inData_202(wire_switch_in_stage5[202]), .inData_203(wire_switch_in_stage5[203]), .inData_204(wire_switch_in_stage5[204]), .inData_205(wire_switch_in_stage5[205]), .inData_206(wire_switch_in_stage5[206]), .inData_207(wire_switch_in_stage5[207]), .inData_208(wire_switch_in_stage5[208]), .inData_209(wire_switch_in_stage5[209]), .inData_210(wire_switch_in_stage5[210]), .inData_211(wire_switch_in_stage5[211]), .inData_212(wire_switch_in_stage5[212]), .inData_213(wire_switch_in_stage5[213]), .inData_214(wire_switch_in_stage5[214]), .inData_215(wire_switch_in_stage5[215]), .inData_216(wire_switch_in_stage5[216]), .inData_217(wire_switch_in_stage5[217]), .inData_218(wire_switch_in_stage5[218]), .inData_219(wire_switch_in_stage5[219]), .inData_220(wire_switch_in_stage5[220]), .inData_221(wire_switch_in_stage5[221]), .inData_222(wire_switch_in_stage5[222]), .inData_223(wire_switch_in_stage5[223]), .inData_224(wire_switch_in_stage5[224]), .inData_225(wire_switch_in_stage5[225]), .inData_226(wire_switch_in_stage5[226]), .inData_227(wire_switch_in_stage5[227]), .inData_228(wire_switch_in_stage5[228]), .inData_229(wire_switch_in_stage5[229]), .inData_230(wire_switch_in_stage5[230]), .inData_231(wire_switch_in_stage5[231]), .inData_232(wire_switch_in_stage5[232]), .inData_233(wire_switch_in_stage5[233]), .inData_234(wire_switch_in_stage5[234]), .inData_235(wire_switch_in_stage5[235]), .inData_236(wire_switch_in_stage5[236]), .inData_237(wire_switch_in_stage5[237]), .inData_238(wire_switch_in_stage5[238]), .inData_239(wire_switch_in_stage5[239]), .inData_240(wire_switch_in_stage5[240]), .inData_241(wire_switch_in_stage5[241]), .inData_242(wire_switch_in_stage5[242]), .inData_243(wire_switch_in_stage5[243]), .inData_244(wire_switch_in_stage5[244]), .inData_245(wire_switch_in_stage5[245]), .inData_246(wire_switch_in_stage5[246]), .inData_247(wire_switch_in_stage5[247]), .inData_248(wire_switch_in_stage5[248]), .inData_249(wire_switch_in_stage5[249]), .inData_250(wire_switch_in_stage5[250]), .inData_251(wire_switch_in_stage5[251]), .inData_252(wire_switch_in_stage5[252]), .inData_253(wire_switch_in_stage5[253]), .inData_254(wire_switch_in_stage5[254]), .inData_255(wire_switch_in_stage5[255]), 
        .outData_0(wire_switch_out_stage5[0]), .outData_1(wire_switch_out_stage5[1]), .outData_2(wire_switch_out_stage5[2]), .outData_3(wire_switch_out_stage5[3]), .outData_4(wire_switch_out_stage5[4]), .outData_5(wire_switch_out_stage5[5]), .outData_6(wire_switch_out_stage5[6]), .outData_7(wire_switch_out_stage5[7]), .outData_8(wire_switch_out_stage5[8]), .outData_9(wire_switch_out_stage5[9]), .outData_10(wire_switch_out_stage5[10]), .outData_11(wire_switch_out_stage5[11]), .outData_12(wire_switch_out_stage5[12]), .outData_13(wire_switch_out_stage5[13]), .outData_14(wire_switch_out_stage5[14]), .outData_15(wire_switch_out_stage5[15]), .outData_16(wire_switch_out_stage5[16]), .outData_17(wire_switch_out_stage5[17]), .outData_18(wire_switch_out_stage5[18]), .outData_19(wire_switch_out_stage5[19]), .outData_20(wire_switch_out_stage5[20]), .outData_21(wire_switch_out_stage5[21]), .outData_22(wire_switch_out_stage5[22]), .outData_23(wire_switch_out_stage5[23]), .outData_24(wire_switch_out_stage5[24]), .outData_25(wire_switch_out_stage5[25]), .outData_26(wire_switch_out_stage5[26]), .outData_27(wire_switch_out_stage5[27]), .outData_28(wire_switch_out_stage5[28]), .outData_29(wire_switch_out_stage5[29]), .outData_30(wire_switch_out_stage5[30]), .outData_31(wire_switch_out_stage5[31]), .outData_32(wire_switch_out_stage5[32]), .outData_33(wire_switch_out_stage5[33]), .outData_34(wire_switch_out_stage5[34]), .outData_35(wire_switch_out_stage5[35]), .outData_36(wire_switch_out_stage5[36]), .outData_37(wire_switch_out_stage5[37]), .outData_38(wire_switch_out_stage5[38]), .outData_39(wire_switch_out_stage5[39]), .outData_40(wire_switch_out_stage5[40]), .outData_41(wire_switch_out_stage5[41]), .outData_42(wire_switch_out_stage5[42]), .outData_43(wire_switch_out_stage5[43]), .outData_44(wire_switch_out_stage5[44]), .outData_45(wire_switch_out_stage5[45]), .outData_46(wire_switch_out_stage5[46]), .outData_47(wire_switch_out_stage5[47]), .outData_48(wire_switch_out_stage5[48]), .outData_49(wire_switch_out_stage5[49]), .outData_50(wire_switch_out_stage5[50]), .outData_51(wire_switch_out_stage5[51]), .outData_52(wire_switch_out_stage5[52]), .outData_53(wire_switch_out_stage5[53]), .outData_54(wire_switch_out_stage5[54]), .outData_55(wire_switch_out_stage5[55]), .outData_56(wire_switch_out_stage5[56]), .outData_57(wire_switch_out_stage5[57]), .outData_58(wire_switch_out_stage5[58]), .outData_59(wire_switch_out_stage5[59]), .outData_60(wire_switch_out_stage5[60]), .outData_61(wire_switch_out_stage5[61]), .outData_62(wire_switch_out_stage5[62]), .outData_63(wire_switch_out_stage5[63]), .outData_64(wire_switch_out_stage5[64]), .outData_65(wire_switch_out_stage5[65]), .outData_66(wire_switch_out_stage5[66]), .outData_67(wire_switch_out_stage5[67]), .outData_68(wire_switch_out_stage5[68]), .outData_69(wire_switch_out_stage5[69]), .outData_70(wire_switch_out_stage5[70]), .outData_71(wire_switch_out_stage5[71]), .outData_72(wire_switch_out_stage5[72]), .outData_73(wire_switch_out_stage5[73]), .outData_74(wire_switch_out_stage5[74]), .outData_75(wire_switch_out_stage5[75]), .outData_76(wire_switch_out_stage5[76]), .outData_77(wire_switch_out_stage5[77]), .outData_78(wire_switch_out_stage5[78]), .outData_79(wire_switch_out_stage5[79]), .outData_80(wire_switch_out_stage5[80]), .outData_81(wire_switch_out_stage5[81]), .outData_82(wire_switch_out_stage5[82]), .outData_83(wire_switch_out_stage5[83]), .outData_84(wire_switch_out_stage5[84]), .outData_85(wire_switch_out_stage5[85]), .outData_86(wire_switch_out_stage5[86]), .outData_87(wire_switch_out_stage5[87]), .outData_88(wire_switch_out_stage5[88]), .outData_89(wire_switch_out_stage5[89]), .outData_90(wire_switch_out_stage5[90]), .outData_91(wire_switch_out_stage5[91]), .outData_92(wire_switch_out_stage5[92]), .outData_93(wire_switch_out_stage5[93]), .outData_94(wire_switch_out_stage5[94]), .outData_95(wire_switch_out_stage5[95]), .outData_96(wire_switch_out_stage5[96]), .outData_97(wire_switch_out_stage5[97]), .outData_98(wire_switch_out_stage5[98]), .outData_99(wire_switch_out_stage5[99]), .outData_100(wire_switch_out_stage5[100]), .outData_101(wire_switch_out_stage5[101]), .outData_102(wire_switch_out_stage5[102]), .outData_103(wire_switch_out_stage5[103]), .outData_104(wire_switch_out_stage5[104]), .outData_105(wire_switch_out_stage5[105]), .outData_106(wire_switch_out_stage5[106]), .outData_107(wire_switch_out_stage5[107]), .outData_108(wire_switch_out_stage5[108]), .outData_109(wire_switch_out_stage5[109]), .outData_110(wire_switch_out_stage5[110]), .outData_111(wire_switch_out_stage5[111]), .outData_112(wire_switch_out_stage5[112]), .outData_113(wire_switch_out_stage5[113]), .outData_114(wire_switch_out_stage5[114]), .outData_115(wire_switch_out_stage5[115]), .outData_116(wire_switch_out_stage5[116]), .outData_117(wire_switch_out_stage5[117]), .outData_118(wire_switch_out_stage5[118]), .outData_119(wire_switch_out_stage5[119]), .outData_120(wire_switch_out_stage5[120]), .outData_121(wire_switch_out_stage5[121]), .outData_122(wire_switch_out_stage5[122]), .outData_123(wire_switch_out_stage5[123]), .outData_124(wire_switch_out_stage5[124]), .outData_125(wire_switch_out_stage5[125]), .outData_126(wire_switch_out_stage5[126]), .outData_127(wire_switch_out_stage5[127]), .outData_128(wire_switch_out_stage5[128]), .outData_129(wire_switch_out_stage5[129]), .outData_130(wire_switch_out_stage5[130]), .outData_131(wire_switch_out_stage5[131]), .outData_132(wire_switch_out_stage5[132]), .outData_133(wire_switch_out_stage5[133]), .outData_134(wire_switch_out_stage5[134]), .outData_135(wire_switch_out_stage5[135]), .outData_136(wire_switch_out_stage5[136]), .outData_137(wire_switch_out_stage5[137]), .outData_138(wire_switch_out_stage5[138]), .outData_139(wire_switch_out_stage5[139]), .outData_140(wire_switch_out_stage5[140]), .outData_141(wire_switch_out_stage5[141]), .outData_142(wire_switch_out_stage5[142]), .outData_143(wire_switch_out_stage5[143]), .outData_144(wire_switch_out_stage5[144]), .outData_145(wire_switch_out_stage5[145]), .outData_146(wire_switch_out_stage5[146]), .outData_147(wire_switch_out_stage5[147]), .outData_148(wire_switch_out_stage5[148]), .outData_149(wire_switch_out_stage5[149]), .outData_150(wire_switch_out_stage5[150]), .outData_151(wire_switch_out_stage5[151]), .outData_152(wire_switch_out_stage5[152]), .outData_153(wire_switch_out_stage5[153]), .outData_154(wire_switch_out_stage5[154]), .outData_155(wire_switch_out_stage5[155]), .outData_156(wire_switch_out_stage5[156]), .outData_157(wire_switch_out_stage5[157]), .outData_158(wire_switch_out_stage5[158]), .outData_159(wire_switch_out_stage5[159]), .outData_160(wire_switch_out_stage5[160]), .outData_161(wire_switch_out_stage5[161]), .outData_162(wire_switch_out_stage5[162]), .outData_163(wire_switch_out_stage5[163]), .outData_164(wire_switch_out_stage5[164]), .outData_165(wire_switch_out_stage5[165]), .outData_166(wire_switch_out_stage5[166]), .outData_167(wire_switch_out_stage5[167]), .outData_168(wire_switch_out_stage5[168]), .outData_169(wire_switch_out_stage5[169]), .outData_170(wire_switch_out_stage5[170]), .outData_171(wire_switch_out_stage5[171]), .outData_172(wire_switch_out_stage5[172]), .outData_173(wire_switch_out_stage5[173]), .outData_174(wire_switch_out_stage5[174]), .outData_175(wire_switch_out_stage5[175]), .outData_176(wire_switch_out_stage5[176]), .outData_177(wire_switch_out_stage5[177]), .outData_178(wire_switch_out_stage5[178]), .outData_179(wire_switch_out_stage5[179]), .outData_180(wire_switch_out_stage5[180]), .outData_181(wire_switch_out_stage5[181]), .outData_182(wire_switch_out_stage5[182]), .outData_183(wire_switch_out_stage5[183]), .outData_184(wire_switch_out_stage5[184]), .outData_185(wire_switch_out_stage5[185]), .outData_186(wire_switch_out_stage5[186]), .outData_187(wire_switch_out_stage5[187]), .outData_188(wire_switch_out_stage5[188]), .outData_189(wire_switch_out_stage5[189]), .outData_190(wire_switch_out_stage5[190]), .outData_191(wire_switch_out_stage5[191]), .outData_192(wire_switch_out_stage5[192]), .outData_193(wire_switch_out_stage5[193]), .outData_194(wire_switch_out_stage5[194]), .outData_195(wire_switch_out_stage5[195]), .outData_196(wire_switch_out_stage5[196]), .outData_197(wire_switch_out_stage5[197]), .outData_198(wire_switch_out_stage5[198]), .outData_199(wire_switch_out_stage5[199]), .outData_200(wire_switch_out_stage5[200]), .outData_201(wire_switch_out_stage5[201]), .outData_202(wire_switch_out_stage5[202]), .outData_203(wire_switch_out_stage5[203]), .outData_204(wire_switch_out_stage5[204]), .outData_205(wire_switch_out_stage5[205]), .outData_206(wire_switch_out_stage5[206]), .outData_207(wire_switch_out_stage5[207]), .outData_208(wire_switch_out_stage5[208]), .outData_209(wire_switch_out_stage5[209]), .outData_210(wire_switch_out_stage5[210]), .outData_211(wire_switch_out_stage5[211]), .outData_212(wire_switch_out_stage5[212]), .outData_213(wire_switch_out_stage5[213]), .outData_214(wire_switch_out_stage5[214]), .outData_215(wire_switch_out_stage5[215]), .outData_216(wire_switch_out_stage5[216]), .outData_217(wire_switch_out_stage5[217]), .outData_218(wire_switch_out_stage5[218]), .outData_219(wire_switch_out_stage5[219]), .outData_220(wire_switch_out_stage5[220]), .outData_221(wire_switch_out_stage5[221]), .outData_222(wire_switch_out_stage5[222]), .outData_223(wire_switch_out_stage5[223]), .outData_224(wire_switch_out_stage5[224]), .outData_225(wire_switch_out_stage5[225]), .outData_226(wire_switch_out_stage5[226]), .outData_227(wire_switch_out_stage5[227]), .outData_228(wire_switch_out_stage5[228]), .outData_229(wire_switch_out_stage5[229]), .outData_230(wire_switch_out_stage5[230]), .outData_231(wire_switch_out_stage5[231]), .outData_232(wire_switch_out_stage5[232]), .outData_233(wire_switch_out_stage5[233]), .outData_234(wire_switch_out_stage5[234]), .outData_235(wire_switch_out_stage5[235]), .outData_236(wire_switch_out_stage5[236]), .outData_237(wire_switch_out_stage5[237]), .outData_238(wire_switch_out_stage5[238]), .outData_239(wire_switch_out_stage5[239]), .outData_240(wire_switch_out_stage5[240]), .outData_241(wire_switch_out_stage5[241]), .outData_242(wire_switch_out_stage5[242]), .outData_243(wire_switch_out_stage5[243]), .outData_244(wire_switch_out_stage5[244]), .outData_245(wire_switch_out_stage5[245]), .outData_246(wire_switch_out_stage5[246]), .outData_247(wire_switch_out_stage5[247]), .outData_248(wire_switch_out_stage5[248]), .outData_249(wire_switch_out_stage5[249]), .outData_250(wire_switch_out_stage5[250]), .outData_251(wire_switch_out_stage5[251]), .outData_252(wire_switch_out_stage5[252]), .outData_253(wire_switch_out_stage5[253]), .outData_254(wire_switch_out_stage5[254]), .outData_255(wire_switch_out_stage5[255]), 
        .in_start(con_in_start_stage5), .out_start(in_start_stage4), .ctrl(wire_ctrl_stage5), .clk(clk), .rst(rst));
  
  wireCon_dp256_st5_R wire_stage_5(
        .inData_0(wire_switch_out_stage6[0]), .inData_1(wire_switch_out_stage6[1]), .inData_2(wire_switch_out_stage6[2]), .inData_3(wire_switch_out_stage6[3]), .inData_4(wire_switch_out_stage6[4]), .inData_5(wire_switch_out_stage6[5]), .inData_6(wire_switch_out_stage6[6]), .inData_7(wire_switch_out_stage6[7]), .inData_8(wire_switch_out_stage6[8]), .inData_9(wire_switch_out_stage6[9]), .inData_10(wire_switch_out_stage6[10]), .inData_11(wire_switch_out_stage6[11]), .inData_12(wire_switch_out_stage6[12]), .inData_13(wire_switch_out_stage6[13]), .inData_14(wire_switch_out_stage6[14]), .inData_15(wire_switch_out_stage6[15]), .inData_16(wire_switch_out_stage6[16]), .inData_17(wire_switch_out_stage6[17]), .inData_18(wire_switch_out_stage6[18]), .inData_19(wire_switch_out_stage6[19]), .inData_20(wire_switch_out_stage6[20]), .inData_21(wire_switch_out_stage6[21]), .inData_22(wire_switch_out_stage6[22]), .inData_23(wire_switch_out_stage6[23]), .inData_24(wire_switch_out_stage6[24]), .inData_25(wire_switch_out_stage6[25]), .inData_26(wire_switch_out_stage6[26]), .inData_27(wire_switch_out_stage6[27]), .inData_28(wire_switch_out_stage6[28]), .inData_29(wire_switch_out_stage6[29]), .inData_30(wire_switch_out_stage6[30]), .inData_31(wire_switch_out_stage6[31]), .inData_32(wire_switch_out_stage6[32]), .inData_33(wire_switch_out_stage6[33]), .inData_34(wire_switch_out_stage6[34]), .inData_35(wire_switch_out_stage6[35]), .inData_36(wire_switch_out_stage6[36]), .inData_37(wire_switch_out_stage6[37]), .inData_38(wire_switch_out_stage6[38]), .inData_39(wire_switch_out_stage6[39]), .inData_40(wire_switch_out_stage6[40]), .inData_41(wire_switch_out_stage6[41]), .inData_42(wire_switch_out_stage6[42]), .inData_43(wire_switch_out_stage6[43]), .inData_44(wire_switch_out_stage6[44]), .inData_45(wire_switch_out_stage6[45]), .inData_46(wire_switch_out_stage6[46]), .inData_47(wire_switch_out_stage6[47]), .inData_48(wire_switch_out_stage6[48]), .inData_49(wire_switch_out_stage6[49]), .inData_50(wire_switch_out_stage6[50]), .inData_51(wire_switch_out_stage6[51]), .inData_52(wire_switch_out_stage6[52]), .inData_53(wire_switch_out_stage6[53]), .inData_54(wire_switch_out_stage6[54]), .inData_55(wire_switch_out_stage6[55]), .inData_56(wire_switch_out_stage6[56]), .inData_57(wire_switch_out_stage6[57]), .inData_58(wire_switch_out_stage6[58]), .inData_59(wire_switch_out_stage6[59]), .inData_60(wire_switch_out_stage6[60]), .inData_61(wire_switch_out_stage6[61]), .inData_62(wire_switch_out_stage6[62]), .inData_63(wire_switch_out_stage6[63]), .inData_64(wire_switch_out_stage6[64]), .inData_65(wire_switch_out_stage6[65]), .inData_66(wire_switch_out_stage6[66]), .inData_67(wire_switch_out_stage6[67]), .inData_68(wire_switch_out_stage6[68]), .inData_69(wire_switch_out_stage6[69]), .inData_70(wire_switch_out_stage6[70]), .inData_71(wire_switch_out_stage6[71]), .inData_72(wire_switch_out_stage6[72]), .inData_73(wire_switch_out_stage6[73]), .inData_74(wire_switch_out_stage6[74]), .inData_75(wire_switch_out_stage6[75]), .inData_76(wire_switch_out_stage6[76]), .inData_77(wire_switch_out_stage6[77]), .inData_78(wire_switch_out_stage6[78]), .inData_79(wire_switch_out_stage6[79]), .inData_80(wire_switch_out_stage6[80]), .inData_81(wire_switch_out_stage6[81]), .inData_82(wire_switch_out_stage6[82]), .inData_83(wire_switch_out_stage6[83]), .inData_84(wire_switch_out_stage6[84]), .inData_85(wire_switch_out_stage6[85]), .inData_86(wire_switch_out_stage6[86]), .inData_87(wire_switch_out_stage6[87]), .inData_88(wire_switch_out_stage6[88]), .inData_89(wire_switch_out_stage6[89]), .inData_90(wire_switch_out_stage6[90]), .inData_91(wire_switch_out_stage6[91]), .inData_92(wire_switch_out_stage6[92]), .inData_93(wire_switch_out_stage6[93]), .inData_94(wire_switch_out_stage6[94]), .inData_95(wire_switch_out_stage6[95]), .inData_96(wire_switch_out_stage6[96]), .inData_97(wire_switch_out_stage6[97]), .inData_98(wire_switch_out_stage6[98]), .inData_99(wire_switch_out_stage6[99]), .inData_100(wire_switch_out_stage6[100]), .inData_101(wire_switch_out_stage6[101]), .inData_102(wire_switch_out_stage6[102]), .inData_103(wire_switch_out_stage6[103]), .inData_104(wire_switch_out_stage6[104]), .inData_105(wire_switch_out_stage6[105]), .inData_106(wire_switch_out_stage6[106]), .inData_107(wire_switch_out_stage6[107]), .inData_108(wire_switch_out_stage6[108]), .inData_109(wire_switch_out_stage6[109]), .inData_110(wire_switch_out_stage6[110]), .inData_111(wire_switch_out_stage6[111]), .inData_112(wire_switch_out_stage6[112]), .inData_113(wire_switch_out_stage6[113]), .inData_114(wire_switch_out_stage6[114]), .inData_115(wire_switch_out_stage6[115]), .inData_116(wire_switch_out_stage6[116]), .inData_117(wire_switch_out_stage6[117]), .inData_118(wire_switch_out_stage6[118]), .inData_119(wire_switch_out_stage6[119]), .inData_120(wire_switch_out_stage6[120]), .inData_121(wire_switch_out_stage6[121]), .inData_122(wire_switch_out_stage6[122]), .inData_123(wire_switch_out_stage6[123]), .inData_124(wire_switch_out_stage6[124]), .inData_125(wire_switch_out_stage6[125]), .inData_126(wire_switch_out_stage6[126]), .inData_127(wire_switch_out_stage6[127]), .inData_128(wire_switch_out_stage6[128]), .inData_129(wire_switch_out_stage6[129]), .inData_130(wire_switch_out_stage6[130]), .inData_131(wire_switch_out_stage6[131]), .inData_132(wire_switch_out_stage6[132]), .inData_133(wire_switch_out_stage6[133]), .inData_134(wire_switch_out_stage6[134]), .inData_135(wire_switch_out_stage6[135]), .inData_136(wire_switch_out_stage6[136]), .inData_137(wire_switch_out_stage6[137]), .inData_138(wire_switch_out_stage6[138]), .inData_139(wire_switch_out_stage6[139]), .inData_140(wire_switch_out_stage6[140]), .inData_141(wire_switch_out_stage6[141]), .inData_142(wire_switch_out_stage6[142]), .inData_143(wire_switch_out_stage6[143]), .inData_144(wire_switch_out_stage6[144]), .inData_145(wire_switch_out_stage6[145]), .inData_146(wire_switch_out_stage6[146]), .inData_147(wire_switch_out_stage6[147]), .inData_148(wire_switch_out_stage6[148]), .inData_149(wire_switch_out_stage6[149]), .inData_150(wire_switch_out_stage6[150]), .inData_151(wire_switch_out_stage6[151]), .inData_152(wire_switch_out_stage6[152]), .inData_153(wire_switch_out_stage6[153]), .inData_154(wire_switch_out_stage6[154]), .inData_155(wire_switch_out_stage6[155]), .inData_156(wire_switch_out_stage6[156]), .inData_157(wire_switch_out_stage6[157]), .inData_158(wire_switch_out_stage6[158]), .inData_159(wire_switch_out_stage6[159]), .inData_160(wire_switch_out_stage6[160]), .inData_161(wire_switch_out_stage6[161]), .inData_162(wire_switch_out_stage6[162]), .inData_163(wire_switch_out_stage6[163]), .inData_164(wire_switch_out_stage6[164]), .inData_165(wire_switch_out_stage6[165]), .inData_166(wire_switch_out_stage6[166]), .inData_167(wire_switch_out_stage6[167]), .inData_168(wire_switch_out_stage6[168]), .inData_169(wire_switch_out_stage6[169]), .inData_170(wire_switch_out_stage6[170]), .inData_171(wire_switch_out_stage6[171]), .inData_172(wire_switch_out_stage6[172]), .inData_173(wire_switch_out_stage6[173]), .inData_174(wire_switch_out_stage6[174]), .inData_175(wire_switch_out_stage6[175]), .inData_176(wire_switch_out_stage6[176]), .inData_177(wire_switch_out_stage6[177]), .inData_178(wire_switch_out_stage6[178]), .inData_179(wire_switch_out_stage6[179]), .inData_180(wire_switch_out_stage6[180]), .inData_181(wire_switch_out_stage6[181]), .inData_182(wire_switch_out_stage6[182]), .inData_183(wire_switch_out_stage6[183]), .inData_184(wire_switch_out_stage6[184]), .inData_185(wire_switch_out_stage6[185]), .inData_186(wire_switch_out_stage6[186]), .inData_187(wire_switch_out_stage6[187]), .inData_188(wire_switch_out_stage6[188]), .inData_189(wire_switch_out_stage6[189]), .inData_190(wire_switch_out_stage6[190]), .inData_191(wire_switch_out_stage6[191]), .inData_192(wire_switch_out_stage6[192]), .inData_193(wire_switch_out_stage6[193]), .inData_194(wire_switch_out_stage6[194]), .inData_195(wire_switch_out_stage6[195]), .inData_196(wire_switch_out_stage6[196]), .inData_197(wire_switch_out_stage6[197]), .inData_198(wire_switch_out_stage6[198]), .inData_199(wire_switch_out_stage6[199]), .inData_200(wire_switch_out_stage6[200]), .inData_201(wire_switch_out_stage6[201]), .inData_202(wire_switch_out_stage6[202]), .inData_203(wire_switch_out_stage6[203]), .inData_204(wire_switch_out_stage6[204]), .inData_205(wire_switch_out_stage6[205]), .inData_206(wire_switch_out_stage6[206]), .inData_207(wire_switch_out_stage6[207]), .inData_208(wire_switch_out_stage6[208]), .inData_209(wire_switch_out_stage6[209]), .inData_210(wire_switch_out_stage6[210]), .inData_211(wire_switch_out_stage6[211]), .inData_212(wire_switch_out_stage6[212]), .inData_213(wire_switch_out_stage6[213]), .inData_214(wire_switch_out_stage6[214]), .inData_215(wire_switch_out_stage6[215]), .inData_216(wire_switch_out_stage6[216]), .inData_217(wire_switch_out_stage6[217]), .inData_218(wire_switch_out_stage6[218]), .inData_219(wire_switch_out_stage6[219]), .inData_220(wire_switch_out_stage6[220]), .inData_221(wire_switch_out_stage6[221]), .inData_222(wire_switch_out_stage6[222]), .inData_223(wire_switch_out_stage6[223]), .inData_224(wire_switch_out_stage6[224]), .inData_225(wire_switch_out_stage6[225]), .inData_226(wire_switch_out_stage6[226]), .inData_227(wire_switch_out_stage6[227]), .inData_228(wire_switch_out_stage6[228]), .inData_229(wire_switch_out_stage6[229]), .inData_230(wire_switch_out_stage6[230]), .inData_231(wire_switch_out_stage6[231]), .inData_232(wire_switch_out_stage6[232]), .inData_233(wire_switch_out_stage6[233]), .inData_234(wire_switch_out_stage6[234]), .inData_235(wire_switch_out_stage6[235]), .inData_236(wire_switch_out_stage6[236]), .inData_237(wire_switch_out_stage6[237]), .inData_238(wire_switch_out_stage6[238]), .inData_239(wire_switch_out_stage6[239]), .inData_240(wire_switch_out_stage6[240]), .inData_241(wire_switch_out_stage6[241]), .inData_242(wire_switch_out_stage6[242]), .inData_243(wire_switch_out_stage6[243]), .inData_244(wire_switch_out_stage6[244]), .inData_245(wire_switch_out_stage6[245]), .inData_246(wire_switch_out_stage6[246]), .inData_247(wire_switch_out_stage6[247]), .inData_248(wire_switch_out_stage6[248]), .inData_249(wire_switch_out_stage6[249]), .inData_250(wire_switch_out_stage6[250]), .inData_251(wire_switch_out_stage6[251]), .inData_252(wire_switch_out_stage6[252]), .inData_253(wire_switch_out_stage6[253]), .inData_254(wire_switch_out_stage6[254]), .inData_255(wire_switch_out_stage6[255]), 
        .outData_0(wire_switch_in_stage5[0]), .outData_1(wire_switch_in_stage5[1]), .outData_2(wire_switch_in_stage5[2]), .outData_3(wire_switch_in_stage5[3]), .outData_4(wire_switch_in_stage5[4]), .outData_5(wire_switch_in_stage5[5]), .outData_6(wire_switch_in_stage5[6]), .outData_7(wire_switch_in_stage5[7]), .outData_8(wire_switch_in_stage5[8]), .outData_9(wire_switch_in_stage5[9]), .outData_10(wire_switch_in_stage5[10]), .outData_11(wire_switch_in_stage5[11]), .outData_12(wire_switch_in_stage5[12]), .outData_13(wire_switch_in_stage5[13]), .outData_14(wire_switch_in_stage5[14]), .outData_15(wire_switch_in_stage5[15]), .outData_16(wire_switch_in_stage5[16]), .outData_17(wire_switch_in_stage5[17]), .outData_18(wire_switch_in_stage5[18]), .outData_19(wire_switch_in_stage5[19]), .outData_20(wire_switch_in_stage5[20]), .outData_21(wire_switch_in_stage5[21]), .outData_22(wire_switch_in_stage5[22]), .outData_23(wire_switch_in_stage5[23]), .outData_24(wire_switch_in_stage5[24]), .outData_25(wire_switch_in_stage5[25]), .outData_26(wire_switch_in_stage5[26]), .outData_27(wire_switch_in_stage5[27]), .outData_28(wire_switch_in_stage5[28]), .outData_29(wire_switch_in_stage5[29]), .outData_30(wire_switch_in_stage5[30]), .outData_31(wire_switch_in_stage5[31]), .outData_32(wire_switch_in_stage5[32]), .outData_33(wire_switch_in_stage5[33]), .outData_34(wire_switch_in_stage5[34]), .outData_35(wire_switch_in_stage5[35]), .outData_36(wire_switch_in_stage5[36]), .outData_37(wire_switch_in_stage5[37]), .outData_38(wire_switch_in_stage5[38]), .outData_39(wire_switch_in_stage5[39]), .outData_40(wire_switch_in_stage5[40]), .outData_41(wire_switch_in_stage5[41]), .outData_42(wire_switch_in_stage5[42]), .outData_43(wire_switch_in_stage5[43]), .outData_44(wire_switch_in_stage5[44]), .outData_45(wire_switch_in_stage5[45]), .outData_46(wire_switch_in_stage5[46]), .outData_47(wire_switch_in_stage5[47]), .outData_48(wire_switch_in_stage5[48]), .outData_49(wire_switch_in_stage5[49]), .outData_50(wire_switch_in_stage5[50]), .outData_51(wire_switch_in_stage5[51]), .outData_52(wire_switch_in_stage5[52]), .outData_53(wire_switch_in_stage5[53]), .outData_54(wire_switch_in_stage5[54]), .outData_55(wire_switch_in_stage5[55]), .outData_56(wire_switch_in_stage5[56]), .outData_57(wire_switch_in_stage5[57]), .outData_58(wire_switch_in_stage5[58]), .outData_59(wire_switch_in_stage5[59]), .outData_60(wire_switch_in_stage5[60]), .outData_61(wire_switch_in_stage5[61]), .outData_62(wire_switch_in_stage5[62]), .outData_63(wire_switch_in_stage5[63]), .outData_64(wire_switch_in_stage5[64]), .outData_65(wire_switch_in_stage5[65]), .outData_66(wire_switch_in_stage5[66]), .outData_67(wire_switch_in_stage5[67]), .outData_68(wire_switch_in_stage5[68]), .outData_69(wire_switch_in_stage5[69]), .outData_70(wire_switch_in_stage5[70]), .outData_71(wire_switch_in_stage5[71]), .outData_72(wire_switch_in_stage5[72]), .outData_73(wire_switch_in_stage5[73]), .outData_74(wire_switch_in_stage5[74]), .outData_75(wire_switch_in_stage5[75]), .outData_76(wire_switch_in_stage5[76]), .outData_77(wire_switch_in_stage5[77]), .outData_78(wire_switch_in_stage5[78]), .outData_79(wire_switch_in_stage5[79]), .outData_80(wire_switch_in_stage5[80]), .outData_81(wire_switch_in_stage5[81]), .outData_82(wire_switch_in_stage5[82]), .outData_83(wire_switch_in_stage5[83]), .outData_84(wire_switch_in_stage5[84]), .outData_85(wire_switch_in_stage5[85]), .outData_86(wire_switch_in_stage5[86]), .outData_87(wire_switch_in_stage5[87]), .outData_88(wire_switch_in_stage5[88]), .outData_89(wire_switch_in_stage5[89]), .outData_90(wire_switch_in_stage5[90]), .outData_91(wire_switch_in_stage5[91]), .outData_92(wire_switch_in_stage5[92]), .outData_93(wire_switch_in_stage5[93]), .outData_94(wire_switch_in_stage5[94]), .outData_95(wire_switch_in_stage5[95]), .outData_96(wire_switch_in_stage5[96]), .outData_97(wire_switch_in_stage5[97]), .outData_98(wire_switch_in_stage5[98]), .outData_99(wire_switch_in_stage5[99]), .outData_100(wire_switch_in_stage5[100]), .outData_101(wire_switch_in_stage5[101]), .outData_102(wire_switch_in_stage5[102]), .outData_103(wire_switch_in_stage5[103]), .outData_104(wire_switch_in_stage5[104]), .outData_105(wire_switch_in_stage5[105]), .outData_106(wire_switch_in_stage5[106]), .outData_107(wire_switch_in_stage5[107]), .outData_108(wire_switch_in_stage5[108]), .outData_109(wire_switch_in_stage5[109]), .outData_110(wire_switch_in_stage5[110]), .outData_111(wire_switch_in_stage5[111]), .outData_112(wire_switch_in_stage5[112]), .outData_113(wire_switch_in_stage5[113]), .outData_114(wire_switch_in_stage5[114]), .outData_115(wire_switch_in_stage5[115]), .outData_116(wire_switch_in_stage5[116]), .outData_117(wire_switch_in_stage5[117]), .outData_118(wire_switch_in_stage5[118]), .outData_119(wire_switch_in_stage5[119]), .outData_120(wire_switch_in_stage5[120]), .outData_121(wire_switch_in_stage5[121]), .outData_122(wire_switch_in_stage5[122]), .outData_123(wire_switch_in_stage5[123]), .outData_124(wire_switch_in_stage5[124]), .outData_125(wire_switch_in_stage5[125]), .outData_126(wire_switch_in_stage5[126]), .outData_127(wire_switch_in_stage5[127]), .outData_128(wire_switch_in_stage5[128]), .outData_129(wire_switch_in_stage5[129]), .outData_130(wire_switch_in_stage5[130]), .outData_131(wire_switch_in_stage5[131]), .outData_132(wire_switch_in_stage5[132]), .outData_133(wire_switch_in_stage5[133]), .outData_134(wire_switch_in_stage5[134]), .outData_135(wire_switch_in_stage5[135]), .outData_136(wire_switch_in_stage5[136]), .outData_137(wire_switch_in_stage5[137]), .outData_138(wire_switch_in_stage5[138]), .outData_139(wire_switch_in_stage5[139]), .outData_140(wire_switch_in_stage5[140]), .outData_141(wire_switch_in_stage5[141]), .outData_142(wire_switch_in_stage5[142]), .outData_143(wire_switch_in_stage5[143]), .outData_144(wire_switch_in_stage5[144]), .outData_145(wire_switch_in_stage5[145]), .outData_146(wire_switch_in_stage5[146]), .outData_147(wire_switch_in_stage5[147]), .outData_148(wire_switch_in_stage5[148]), .outData_149(wire_switch_in_stage5[149]), .outData_150(wire_switch_in_stage5[150]), .outData_151(wire_switch_in_stage5[151]), .outData_152(wire_switch_in_stage5[152]), .outData_153(wire_switch_in_stage5[153]), .outData_154(wire_switch_in_stage5[154]), .outData_155(wire_switch_in_stage5[155]), .outData_156(wire_switch_in_stage5[156]), .outData_157(wire_switch_in_stage5[157]), .outData_158(wire_switch_in_stage5[158]), .outData_159(wire_switch_in_stage5[159]), .outData_160(wire_switch_in_stage5[160]), .outData_161(wire_switch_in_stage5[161]), .outData_162(wire_switch_in_stage5[162]), .outData_163(wire_switch_in_stage5[163]), .outData_164(wire_switch_in_stage5[164]), .outData_165(wire_switch_in_stage5[165]), .outData_166(wire_switch_in_stage5[166]), .outData_167(wire_switch_in_stage5[167]), .outData_168(wire_switch_in_stage5[168]), .outData_169(wire_switch_in_stage5[169]), .outData_170(wire_switch_in_stage5[170]), .outData_171(wire_switch_in_stage5[171]), .outData_172(wire_switch_in_stage5[172]), .outData_173(wire_switch_in_stage5[173]), .outData_174(wire_switch_in_stage5[174]), .outData_175(wire_switch_in_stage5[175]), .outData_176(wire_switch_in_stage5[176]), .outData_177(wire_switch_in_stage5[177]), .outData_178(wire_switch_in_stage5[178]), .outData_179(wire_switch_in_stage5[179]), .outData_180(wire_switch_in_stage5[180]), .outData_181(wire_switch_in_stage5[181]), .outData_182(wire_switch_in_stage5[182]), .outData_183(wire_switch_in_stage5[183]), .outData_184(wire_switch_in_stage5[184]), .outData_185(wire_switch_in_stage5[185]), .outData_186(wire_switch_in_stage5[186]), .outData_187(wire_switch_in_stage5[187]), .outData_188(wire_switch_in_stage5[188]), .outData_189(wire_switch_in_stage5[189]), .outData_190(wire_switch_in_stage5[190]), .outData_191(wire_switch_in_stage5[191]), .outData_192(wire_switch_in_stage5[192]), .outData_193(wire_switch_in_stage5[193]), .outData_194(wire_switch_in_stage5[194]), .outData_195(wire_switch_in_stage5[195]), .outData_196(wire_switch_in_stage5[196]), .outData_197(wire_switch_in_stage5[197]), .outData_198(wire_switch_in_stage5[198]), .outData_199(wire_switch_in_stage5[199]), .outData_200(wire_switch_in_stage5[200]), .outData_201(wire_switch_in_stage5[201]), .outData_202(wire_switch_in_stage5[202]), .outData_203(wire_switch_in_stage5[203]), .outData_204(wire_switch_in_stage5[204]), .outData_205(wire_switch_in_stage5[205]), .outData_206(wire_switch_in_stage5[206]), .outData_207(wire_switch_in_stage5[207]), .outData_208(wire_switch_in_stage5[208]), .outData_209(wire_switch_in_stage5[209]), .outData_210(wire_switch_in_stage5[210]), .outData_211(wire_switch_in_stage5[211]), .outData_212(wire_switch_in_stage5[212]), .outData_213(wire_switch_in_stage5[213]), .outData_214(wire_switch_in_stage5[214]), .outData_215(wire_switch_in_stage5[215]), .outData_216(wire_switch_in_stage5[216]), .outData_217(wire_switch_in_stage5[217]), .outData_218(wire_switch_in_stage5[218]), .outData_219(wire_switch_in_stage5[219]), .outData_220(wire_switch_in_stage5[220]), .outData_221(wire_switch_in_stage5[221]), .outData_222(wire_switch_in_stage5[222]), .outData_223(wire_switch_in_stage5[223]), .outData_224(wire_switch_in_stage5[224]), .outData_225(wire_switch_in_stage5[225]), .outData_226(wire_switch_in_stage5[226]), .outData_227(wire_switch_in_stage5[227]), .outData_228(wire_switch_in_stage5[228]), .outData_229(wire_switch_in_stage5[229]), .outData_230(wire_switch_in_stage5[230]), .outData_231(wire_switch_in_stage5[231]), .outData_232(wire_switch_in_stage5[232]), .outData_233(wire_switch_in_stage5[233]), .outData_234(wire_switch_in_stage5[234]), .outData_235(wire_switch_in_stage5[235]), .outData_236(wire_switch_in_stage5[236]), .outData_237(wire_switch_in_stage5[237]), .outData_238(wire_switch_in_stage5[238]), .outData_239(wire_switch_in_stage5[239]), .outData_240(wire_switch_in_stage5[240]), .outData_241(wire_switch_in_stage5[241]), .outData_242(wire_switch_in_stage5[242]), .outData_243(wire_switch_in_stage5[243]), .outData_244(wire_switch_in_stage5[244]), .outData_245(wire_switch_in_stage5[245]), .outData_246(wire_switch_in_stage5[246]), .outData_247(wire_switch_in_stage5[247]), .outData_248(wire_switch_in_stage5[248]), .outData_249(wire_switch_in_stage5[249]), .outData_250(wire_switch_in_stage5[250]), .outData_251(wire_switch_in_stage5[251]), .outData_252(wire_switch_in_stage5[252]), .outData_253(wire_switch_in_stage5[253]), .outData_254(wire_switch_in_stage5[254]), .outData_255(wire_switch_in_stage5[255]), 
        .in_start(in_start_stage5), .out_start(con_in_start_stage5), .clk(clk), .rst(rst)); 

  
  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[0] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[1] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[2] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[3] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[4] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[5] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[6] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[7] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[8] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[9] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[10] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[11] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[12] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[13] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[14] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[15] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[16] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[17] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[18] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[19] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[20] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[21] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[22] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[23] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[24] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[25] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[26] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[27] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[28] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[29] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[30] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[31] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[32] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[33] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[34] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[35] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[36] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[37] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[38] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[39] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[40] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[41] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[42] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[43] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[44] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[45] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[46] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[47] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[48] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[49] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[50] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[51] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[52] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[53] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[54] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[55] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[56] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[57] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[58] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[59] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[60] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[61] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[62] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[63] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[64] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[65] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[66] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[67] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[68] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[69] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[70] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[71] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[72] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[73] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[74] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[75] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[76] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[77] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[78] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[79] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[80] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[81] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[82] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[83] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[84] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[85] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[86] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[87] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[88] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[89] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[90] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[91] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[92] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[93] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[94] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[95] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[96] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[97] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[98] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[99] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[100] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[101] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[102] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[103] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[104] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[105] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[106] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[107] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[108] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[109] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[110] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[111] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[112] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[113] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[114] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[115] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[116] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[117] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[118] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[119] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[120] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[121] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[122] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[123] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[124] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[125] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[126] <= counter_w[2]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage5[127] <= counter_w[2]; 
  end                            

  wire [DATA_WIDTH-1:0] wire_switch_in_stage4[255:0];
  wire [DATA_WIDTH-1:0] wire_switch_out_stage4[255:0];
  reg [127:0] wire_ctrl_stage4;

  switches_stage_st4_0_R switch_stage_4(
        .inData_0(wire_switch_in_stage4[0]), .inData_1(wire_switch_in_stage4[1]), .inData_2(wire_switch_in_stage4[2]), .inData_3(wire_switch_in_stage4[3]), .inData_4(wire_switch_in_stage4[4]), .inData_5(wire_switch_in_stage4[5]), .inData_6(wire_switch_in_stage4[6]), .inData_7(wire_switch_in_stage4[7]), .inData_8(wire_switch_in_stage4[8]), .inData_9(wire_switch_in_stage4[9]), .inData_10(wire_switch_in_stage4[10]), .inData_11(wire_switch_in_stage4[11]), .inData_12(wire_switch_in_stage4[12]), .inData_13(wire_switch_in_stage4[13]), .inData_14(wire_switch_in_stage4[14]), .inData_15(wire_switch_in_stage4[15]), .inData_16(wire_switch_in_stage4[16]), .inData_17(wire_switch_in_stage4[17]), .inData_18(wire_switch_in_stage4[18]), .inData_19(wire_switch_in_stage4[19]), .inData_20(wire_switch_in_stage4[20]), .inData_21(wire_switch_in_stage4[21]), .inData_22(wire_switch_in_stage4[22]), .inData_23(wire_switch_in_stage4[23]), .inData_24(wire_switch_in_stage4[24]), .inData_25(wire_switch_in_stage4[25]), .inData_26(wire_switch_in_stage4[26]), .inData_27(wire_switch_in_stage4[27]), .inData_28(wire_switch_in_stage4[28]), .inData_29(wire_switch_in_stage4[29]), .inData_30(wire_switch_in_stage4[30]), .inData_31(wire_switch_in_stage4[31]), .inData_32(wire_switch_in_stage4[32]), .inData_33(wire_switch_in_stage4[33]), .inData_34(wire_switch_in_stage4[34]), .inData_35(wire_switch_in_stage4[35]), .inData_36(wire_switch_in_stage4[36]), .inData_37(wire_switch_in_stage4[37]), .inData_38(wire_switch_in_stage4[38]), .inData_39(wire_switch_in_stage4[39]), .inData_40(wire_switch_in_stage4[40]), .inData_41(wire_switch_in_stage4[41]), .inData_42(wire_switch_in_stage4[42]), .inData_43(wire_switch_in_stage4[43]), .inData_44(wire_switch_in_stage4[44]), .inData_45(wire_switch_in_stage4[45]), .inData_46(wire_switch_in_stage4[46]), .inData_47(wire_switch_in_stage4[47]), .inData_48(wire_switch_in_stage4[48]), .inData_49(wire_switch_in_stage4[49]), .inData_50(wire_switch_in_stage4[50]), .inData_51(wire_switch_in_stage4[51]), .inData_52(wire_switch_in_stage4[52]), .inData_53(wire_switch_in_stage4[53]), .inData_54(wire_switch_in_stage4[54]), .inData_55(wire_switch_in_stage4[55]), .inData_56(wire_switch_in_stage4[56]), .inData_57(wire_switch_in_stage4[57]), .inData_58(wire_switch_in_stage4[58]), .inData_59(wire_switch_in_stage4[59]), .inData_60(wire_switch_in_stage4[60]), .inData_61(wire_switch_in_stage4[61]), .inData_62(wire_switch_in_stage4[62]), .inData_63(wire_switch_in_stage4[63]), .inData_64(wire_switch_in_stage4[64]), .inData_65(wire_switch_in_stage4[65]), .inData_66(wire_switch_in_stage4[66]), .inData_67(wire_switch_in_stage4[67]), .inData_68(wire_switch_in_stage4[68]), .inData_69(wire_switch_in_stage4[69]), .inData_70(wire_switch_in_stage4[70]), .inData_71(wire_switch_in_stage4[71]), .inData_72(wire_switch_in_stage4[72]), .inData_73(wire_switch_in_stage4[73]), .inData_74(wire_switch_in_stage4[74]), .inData_75(wire_switch_in_stage4[75]), .inData_76(wire_switch_in_stage4[76]), .inData_77(wire_switch_in_stage4[77]), .inData_78(wire_switch_in_stage4[78]), .inData_79(wire_switch_in_stage4[79]), .inData_80(wire_switch_in_stage4[80]), .inData_81(wire_switch_in_stage4[81]), .inData_82(wire_switch_in_stage4[82]), .inData_83(wire_switch_in_stage4[83]), .inData_84(wire_switch_in_stage4[84]), .inData_85(wire_switch_in_stage4[85]), .inData_86(wire_switch_in_stage4[86]), .inData_87(wire_switch_in_stage4[87]), .inData_88(wire_switch_in_stage4[88]), .inData_89(wire_switch_in_stage4[89]), .inData_90(wire_switch_in_stage4[90]), .inData_91(wire_switch_in_stage4[91]), .inData_92(wire_switch_in_stage4[92]), .inData_93(wire_switch_in_stage4[93]), .inData_94(wire_switch_in_stage4[94]), .inData_95(wire_switch_in_stage4[95]), .inData_96(wire_switch_in_stage4[96]), .inData_97(wire_switch_in_stage4[97]), .inData_98(wire_switch_in_stage4[98]), .inData_99(wire_switch_in_stage4[99]), .inData_100(wire_switch_in_stage4[100]), .inData_101(wire_switch_in_stage4[101]), .inData_102(wire_switch_in_stage4[102]), .inData_103(wire_switch_in_stage4[103]), .inData_104(wire_switch_in_stage4[104]), .inData_105(wire_switch_in_stage4[105]), .inData_106(wire_switch_in_stage4[106]), .inData_107(wire_switch_in_stage4[107]), .inData_108(wire_switch_in_stage4[108]), .inData_109(wire_switch_in_stage4[109]), .inData_110(wire_switch_in_stage4[110]), .inData_111(wire_switch_in_stage4[111]), .inData_112(wire_switch_in_stage4[112]), .inData_113(wire_switch_in_stage4[113]), .inData_114(wire_switch_in_stage4[114]), .inData_115(wire_switch_in_stage4[115]), .inData_116(wire_switch_in_stage4[116]), .inData_117(wire_switch_in_stage4[117]), .inData_118(wire_switch_in_stage4[118]), .inData_119(wire_switch_in_stage4[119]), .inData_120(wire_switch_in_stage4[120]), .inData_121(wire_switch_in_stage4[121]), .inData_122(wire_switch_in_stage4[122]), .inData_123(wire_switch_in_stage4[123]), .inData_124(wire_switch_in_stage4[124]), .inData_125(wire_switch_in_stage4[125]), .inData_126(wire_switch_in_stage4[126]), .inData_127(wire_switch_in_stage4[127]), .inData_128(wire_switch_in_stage4[128]), .inData_129(wire_switch_in_stage4[129]), .inData_130(wire_switch_in_stage4[130]), .inData_131(wire_switch_in_stage4[131]), .inData_132(wire_switch_in_stage4[132]), .inData_133(wire_switch_in_stage4[133]), .inData_134(wire_switch_in_stage4[134]), .inData_135(wire_switch_in_stage4[135]), .inData_136(wire_switch_in_stage4[136]), .inData_137(wire_switch_in_stage4[137]), .inData_138(wire_switch_in_stage4[138]), .inData_139(wire_switch_in_stage4[139]), .inData_140(wire_switch_in_stage4[140]), .inData_141(wire_switch_in_stage4[141]), .inData_142(wire_switch_in_stage4[142]), .inData_143(wire_switch_in_stage4[143]), .inData_144(wire_switch_in_stage4[144]), .inData_145(wire_switch_in_stage4[145]), .inData_146(wire_switch_in_stage4[146]), .inData_147(wire_switch_in_stage4[147]), .inData_148(wire_switch_in_stage4[148]), .inData_149(wire_switch_in_stage4[149]), .inData_150(wire_switch_in_stage4[150]), .inData_151(wire_switch_in_stage4[151]), .inData_152(wire_switch_in_stage4[152]), .inData_153(wire_switch_in_stage4[153]), .inData_154(wire_switch_in_stage4[154]), .inData_155(wire_switch_in_stage4[155]), .inData_156(wire_switch_in_stage4[156]), .inData_157(wire_switch_in_stage4[157]), .inData_158(wire_switch_in_stage4[158]), .inData_159(wire_switch_in_stage4[159]), .inData_160(wire_switch_in_stage4[160]), .inData_161(wire_switch_in_stage4[161]), .inData_162(wire_switch_in_stage4[162]), .inData_163(wire_switch_in_stage4[163]), .inData_164(wire_switch_in_stage4[164]), .inData_165(wire_switch_in_stage4[165]), .inData_166(wire_switch_in_stage4[166]), .inData_167(wire_switch_in_stage4[167]), .inData_168(wire_switch_in_stage4[168]), .inData_169(wire_switch_in_stage4[169]), .inData_170(wire_switch_in_stage4[170]), .inData_171(wire_switch_in_stage4[171]), .inData_172(wire_switch_in_stage4[172]), .inData_173(wire_switch_in_stage4[173]), .inData_174(wire_switch_in_stage4[174]), .inData_175(wire_switch_in_stage4[175]), .inData_176(wire_switch_in_stage4[176]), .inData_177(wire_switch_in_stage4[177]), .inData_178(wire_switch_in_stage4[178]), .inData_179(wire_switch_in_stage4[179]), .inData_180(wire_switch_in_stage4[180]), .inData_181(wire_switch_in_stage4[181]), .inData_182(wire_switch_in_stage4[182]), .inData_183(wire_switch_in_stage4[183]), .inData_184(wire_switch_in_stage4[184]), .inData_185(wire_switch_in_stage4[185]), .inData_186(wire_switch_in_stage4[186]), .inData_187(wire_switch_in_stage4[187]), .inData_188(wire_switch_in_stage4[188]), .inData_189(wire_switch_in_stage4[189]), .inData_190(wire_switch_in_stage4[190]), .inData_191(wire_switch_in_stage4[191]), .inData_192(wire_switch_in_stage4[192]), .inData_193(wire_switch_in_stage4[193]), .inData_194(wire_switch_in_stage4[194]), .inData_195(wire_switch_in_stage4[195]), .inData_196(wire_switch_in_stage4[196]), .inData_197(wire_switch_in_stage4[197]), .inData_198(wire_switch_in_stage4[198]), .inData_199(wire_switch_in_stage4[199]), .inData_200(wire_switch_in_stage4[200]), .inData_201(wire_switch_in_stage4[201]), .inData_202(wire_switch_in_stage4[202]), .inData_203(wire_switch_in_stage4[203]), .inData_204(wire_switch_in_stage4[204]), .inData_205(wire_switch_in_stage4[205]), .inData_206(wire_switch_in_stage4[206]), .inData_207(wire_switch_in_stage4[207]), .inData_208(wire_switch_in_stage4[208]), .inData_209(wire_switch_in_stage4[209]), .inData_210(wire_switch_in_stage4[210]), .inData_211(wire_switch_in_stage4[211]), .inData_212(wire_switch_in_stage4[212]), .inData_213(wire_switch_in_stage4[213]), .inData_214(wire_switch_in_stage4[214]), .inData_215(wire_switch_in_stage4[215]), .inData_216(wire_switch_in_stage4[216]), .inData_217(wire_switch_in_stage4[217]), .inData_218(wire_switch_in_stage4[218]), .inData_219(wire_switch_in_stage4[219]), .inData_220(wire_switch_in_stage4[220]), .inData_221(wire_switch_in_stage4[221]), .inData_222(wire_switch_in_stage4[222]), .inData_223(wire_switch_in_stage4[223]), .inData_224(wire_switch_in_stage4[224]), .inData_225(wire_switch_in_stage4[225]), .inData_226(wire_switch_in_stage4[226]), .inData_227(wire_switch_in_stage4[227]), .inData_228(wire_switch_in_stage4[228]), .inData_229(wire_switch_in_stage4[229]), .inData_230(wire_switch_in_stage4[230]), .inData_231(wire_switch_in_stage4[231]), .inData_232(wire_switch_in_stage4[232]), .inData_233(wire_switch_in_stage4[233]), .inData_234(wire_switch_in_stage4[234]), .inData_235(wire_switch_in_stage4[235]), .inData_236(wire_switch_in_stage4[236]), .inData_237(wire_switch_in_stage4[237]), .inData_238(wire_switch_in_stage4[238]), .inData_239(wire_switch_in_stage4[239]), .inData_240(wire_switch_in_stage4[240]), .inData_241(wire_switch_in_stage4[241]), .inData_242(wire_switch_in_stage4[242]), .inData_243(wire_switch_in_stage4[243]), .inData_244(wire_switch_in_stage4[244]), .inData_245(wire_switch_in_stage4[245]), .inData_246(wire_switch_in_stage4[246]), .inData_247(wire_switch_in_stage4[247]), .inData_248(wire_switch_in_stage4[248]), .inData_249(wire_switch_in_stage4[249]), .inData_250(wire_switch_in_stage4[250]), .inData_251(wire_switch_in_stage4[251]), .inData_252(wire_switch_in_stage4[252]), .inData_253(wire_switch_in_stage4[253]), .inData_254(wire_switch_in_stage4[254]), .inData_255(wire_switch_in_stage4[255]), 
        .outData_0(wire_switch_out_stage4[0]), .outData_1(wire_switch_out_stage4[1]), .outData_2(wire_switch_out_stage4[2]), .outData_3(wire_switch_out_stage4[3]), .outData_4(wire_switch_out_stage4[4]), .outData_5(wire_switch_out_stage4[5]), .outData_6(wire_switch_out_stage4[6]), .outData_7(wire_switch_out_stage4[7]), .outData_8(wire_switch_out_stage4[8]), .outData_9(wire_switch_out_stage4[9]), .outData_10(wire_switch_out_stage4[10]), .outData_11(wire_switch_out_stage4[11]), .outData_12(wire_switch_out_stage4[12]), .outData_13(wire_switch_out_stage4[13]), .outData_14(wire_switch_out_stage4[14]), .outData_15(wire_switch_out_stage4[15]), .outData_16(wire_switch_out_stage4[16]), .outData_17(wire_switch_out_stage4[17]), .outData_18(wire_switch_out_stage4[18]), .outData_19(wire_switch_out_stage4[19]), .outData_20(wire_switch_out_stage4[20]), .outData_21(wire_switch_out_stage4[21]), .outData_22(wire_switch_out_stage4[22]), .outData_23(wire_switch_out_stage4[23]), .outData_24(wire_switch_out_stage4[24]), .outData_25(wire_switch_out_stage4[25]), .outData_26(wire_switch_out_stage4[26]), .outData_27(wire_switch_out_stage4[27]), .outData_28(wire_switch_out_stage4[28]), .outData_29(wire_switch_out_stage4[29]), .outData_30(wire_switch_out_stage4[30]), .outData_31(wire_switch_out_stage4[31]), .outData_32(wire_switch_out_stage4[32]), .outData_33(wire_switch_out_stage4[33]), .outData_34(wire_switch_out_stage4[34]), .outData_35(wire_switch_out_stage4[35]), .outData_36(wire_switch_out_stage4[36]), .outData_37(wire_switch_out_stage4[37]), .outData_38(wire_switch_out_stage4[38]), .outData_39(wire_switch_out_stage4[39]), .outData_40(wire_switch_out_stage4[40]), .outData_41(wire_switch_out_stage4[41]), .outData_42(wire_switch_out_stage4[42]), .outData_43(wire_switch_out_stage4[43]), .outData_44(wire_switch_out_stage4[44]), .outData_45(wire_switch_out_stage4[45]), .outData_46(wire_switch_out_stage4[46]), .outData_47(wire_switch_out_stage4[47]), .outData_48(wire_switch_out_stage4[48]), .outData_49(wire_switch_out_stage4[49]), .outData_50(wire_switch_out_stage4[50]), .outData_51(wire_switch_out_stage4[51]), .outData_52(wire_switch_out_stage4[52]), .outData_53(wire_switch_out_stage4[53]), .outData_54(wire_switch_out_stage4[54]), .outData_55(wire_switch_out_stage4[55]), .outData_56(wire_switch_out_stage4[56]), .outData_57(wire_switch_out_stage4[57]), .outData_58(wire_switch_out_stage4[58]), .outData_59(wire_switch_out_stage4[59]), .outData_60(wire_switch_out_stage4[60]), .outData_61(wire_switch_out_stage4[61]), .outData_62(wire_switch_out_stage4[62]), .outData_63(wire_switch_out_stage4[63]), .outData_64(wire_switch_out_stage4[64]), .outData_65(wire_switch_out_stage4[65]), .outData_66(wire_switch_out_stage4[66]), .outData_67(wire_switch_out_stage4[67]), .outData_68(wire_switch_out_stage4[68]), .outData_69(wire_switch_out_stage4[69]), .outData_70(wire_switch_out_stage4[70]), .outData_71(wire_switch_out_stage4[71]), .outData_72(wire_switch_out_stage4[72]), .outData_73(wire_switch_out_stage4[73]), .outData_74(wire_switch_out_stage4[74]), .outData_75(wire_switch_out_stage4[75]), .outData_76(wire_switch_out_stage4[76]), .outData_77(wire_switch_out_stage4[77]), .outData_78(wire_switch_out_stage4[78]), .outData_79(wire_switch_out_stage4[79]), .outData_80(wire_switch_out_stage4[80]), .outData_81(wire_switch_out_stage4[81]), .outData_82(wire_switch_out_stage4[82]), .outData_83(wire_switch_out_stage4[83]), .outData_84(wire_switch_out_stage4[84]), .outData_85(wire_switch_out_stage4[85]), .outData_86(wire_switch_out_stage4[86]), .outData_87(wire_switch_out_stage4[87]), .outData_88(wire_switch_out_stage4[88]), .outData_89(wire_switch_out_stage4[89]), .outData_90(wire_switch_out_stage4[90]), .outData_91(wire_switch_out_stage4[91]), .outData_92(wire_switch_out_stage4[92]), .outData_93(wire_switch_out_stage4[93]), .outData_94(wire_switch_out_stage4[94]), .outData_95(wire_switch_out_stage4[95]), .outData_96(wire_switch_out_stage4[96]), .outData_97(wire_switch_out_stage4[97]), .outData_98(wire_switch_out_stage4[98]), .outData_99(wire_switch_out_stage4[99]), .outData_100(wire_switch_out_stage4[100]), .outData_101(wire_switch_out_stage4[101]), .outData_102(wire_switch_out_stage4[102]), .outData_103(wire_switch_out_stage4[103]), .outData_104(wire_switch_out_stage4[104]), .outData_105(wire_switch_out_stage4[105]), .outData_106(wire_switch_out_stage4[106]), .outData_107(wire_switch_out_stage4[107]), .outData_108(wire_switch_out_stage4[108]), .outData_109(wire_switch_out_stage4[109]), .outData_110(wire_switch_out_stage4[110]), .outData_111(wire_switch_out_stage4[111]), .outData_112(wire_switch_out_stage4[112]), .outData_113(wire_switch_out_stage4[113]), .outData_114(wire_switch_out_stage4[114]), .outData_115(wire_switch_out_stage4[115]), .outData_116(wire_switch_out_stage4[116]), .outData_117(wire_switch_out_stage4[117]), .outData_118(wire_switch_out_stage4[118]), .outData_119(wire_switch_out_stage4[119]), .outData_120(wire_switch_out_stage4[120]), .outData_121(wire_switch_out_stage4[121]), .outData_122(wire_switch_out_stage4[122]), .outData_123(wire_switch_out_stage4[123]), .outData_124(wire_switch_out_stage4[124]), .outData_125(wire_switch_out_stage4[125]), .outData_126(wire_switch_out_stage4[126]), .outData_127(wire_switch_out_stage4[127]), .outData_128(wire_switch_out_stage4[128]), .outData_129(wire_switch_out_stage4[129]), .outData_130(wire_switch_out_stage4[130]), .outData_131(wire_switch_out_stage4[131]), .outData_132(wire_switch_out_stage4[132]), .outData_133(wire_switch_out_stage4[133]), .outData_134(wire_switch_out_stage4[134]), .outData_135(wire_switch_out_stage4[135]), .outData_136(wire_switch_out_stage4[136]), .outData_137(wire_switch_out_stage4[137]), .outData_138(wire_switch_out_stage4[138]), .outData_139(wire_switch_out_stage4[139]), .outData_140(wire_switch_out_stage4[140]), .outData_141(wire_switch_out_stage4[141]), .outData_142(wire_switch_out_stage4[142]), .outData_143(wire_switch_out_stage4[143]), .outData_144(wire_switch_out_stage4[144]), .outData_145(wire_switch_out_stage4[145]), .outData_146(wire_switch_out_stage4[146]), .outData_147(wire_switch_out_stage4[147]), .outData_148(wire_switch_out_stage4[148]), .outData_149(wire_switch_out_stage4[149]), .outData_150(wire_switch_out_stage4[150]), .outData_151(wire_switch_out_stage4[151]), .outData_152(wire_switch_out_stage4[152]), .outData_153(wire_switch_out_stage4[153]), .outData_154(wire_switch_out_stage4[154]), .outData_155(wire_switch_out_stage4[155]), .outData_156(wire_switch_out_stage4[156]), .outData_157(wire_switch_out_stage4[157]), .outData_158(wire_switch_out_stage4[158]), .outData_159(wire_switch_out_stage4[159]), .outData_160(wire_switch_out_stage4[160]), .outData_161(wire_switch_out_stage4[161]), .outData_162(wire_switch_out_stage4[162]), .outData_163(wire_switch_out_stage4[163]), .outData_164(wire_switch_out_stage4[164]), .outData_165(wire_switch_out_stage4[165]), .outData_166(wire_switch_out_stage4[166]), .outData_167(wire_switch_out_stage4[167]), .outData_168(wire_switch_out_stage4[168]), .outData_169(wire_switch_out_stage4[169]), .outData_170(wire_switch_out_stage4[170]), .outData_171(wire_switch_out_stage4[171]), .outData_172(wire_switch_out_stage4[172]), .outData_173(wire_switch_out_stage4[173]), .outData_174(wire_switch_out_stage4[174]), .outData_175(wire_switch_out_stage4[175]), .outData_176(wire_switch_out_stage4[176]), .outData_177(wire_switch_out_stage4[177]), .outData_178(wire_switch_out_stage4[178]), .outData_179(wire_switch_out_stage4[179]), .outData_180(wire_switch_out_stage4[180]), .outData_181(wire_switch_out_stage4[181]), .outData_182(wire_switch_out_stage4[182]), .outData_183(wire_switch_out_stage4[183]), .outData_184(wire_switch_out_stage4[184]), .outData_185(wire_switch_out_stage4[185]), .outData_186(wire_switch_out_stage4[186]), .outData_187(wire_switch_out_stage4[187]), .outData_188(wire_switch_out_stage4[188]), .outData_189(wire_switch_out_stage4[189]), .outData_190(wire_switch_out_stage4[190]), .outData_191(wire_switch_out_stage4[191]), .outData_192(wire_switch_out_stage4[192]), .outData_193(wire_switch_out_stage4[193]), .outData_194(wire_switch_out_stage4[194]), .outData_195(wire_switch_out_stage4[195]), .outData_196(wire_switch_out_stage4[196]), .outData_197(wire_switch_out_stage4[197]), .outData_198(wire_switch_out_stage4[198]), .outData_199(wire_switch_out_stage4[199]), .outData_200(wire_switch_out_stage4[200]), .outData_201(wire_switch_out_stage4[201]), .outData_202(wire_switch_out_stage4[202]), .outData_203(wire_switch_out_stage4[203]), .outData_204(wire_switch_out_stage4[204]), .outData_205(wire_switch_out_stage4[205]), .outData_206(wire_switch_out_stage4[206]), .outData_207(wire_switch_out_stage4[207]), .outData_208(wire_switch_out_stage4[208]), .outData_209(wire_switch_out_stage4[209]), .outData_210(wire_switch_out_stage4[210]), .outData_211(wire_switch_out_stage4[211]), .outData_212(wire_switch_out_stage4[212]), .outData_213(wire_switch_out_stage4[213]), .outData_214(wire_switch_out_stage4[214]), .outData_215(wire_switch_out_stage4[215]), .outData_216(wire_switch_out_stage4[216]), .outData_217(wire_switch_out_stage4[217]), .outData_218(wire_switch_out_stage4[218]), .outData_219(wire_switch_out_stage4[219]), .outData_220(wire_switch_out_stage4[220]), .outData_221(wire_switch_out_stage4[221]), .outData_222(wire_switch_out_stage4[222]), .outData_223(wire_switch_out_stage4[223]), .outData_224(wire_switch_out_stage4[224]), .outData_225(wire_switch_out_stage4[225]), .outData_226(wire_switch_out_stage4[226]), .outData_227(wire_switch_out_stage4[227]), .outData_228(wire_switch_out_stage4[228]), .outData_229(wire_switch_out_stage4[229]), .outData_230(wire_switch_out_stage4[230]), .outData_231(wire_switch_out_stage4[231]), .outData_232(wire_switch_out_stage4[232]), .outData_233(wire_switch_out_stage4[233]), .outData_234(wire_switch_out_stage4[234]), .outData_235(wire_switch_out_stage4[235]), .outData_236(wire_switch_out_stage4[236]), .outData_237(wire_switch_out_stage4[237]), .outData_238(wire_switch_out_stage4[238]), .outData_239(wire_switch_out_stage4[239]), .outData_240(wire_switch_out_stage4[240]), .outData_241(wire_switch_out_stage4[241]), .outData_242(wire_switch_out_stage4[242]), .outData_243(wire_switch_out_stage4[243]), .outData_244(wire_switch_out_stage4[244]), .outData_245(wire_switch_out_stage4[245]), .outData_246(wire_switch_out_stage4[246]), .outData_247(wire_switch_out_stage4[247]), .outData_248(wire_switch_out_stage4[248]), .outData_249(wire_switch_out_stage4[249]), .outData_250(wire_switch_out_stage4[250]), .outData_251(wire_switch_out_stage4[251]), .outData_252(wire_switch_out_stage4[252]), .outData_253(wire_switch_out_stage4[253]), .outData_254(wire_switch_out_stage4[254]), .outData_255(wire_switch_out_stage4[255]), 
        .in_start(con_in_start_stage4), .out_start(in_start_stage3), .ctrl(wire_ctrl_stage4), .clk(clk), .rst(rst));
  
  wireCon_dp256_st4_R wire_stage_4(
        .inData_0(wire_switch_out_stage5[0]), .inData_1(wire_switch_out_stage5[1]), .inData_2(wire_switch_out_stage5[2]), .inData_3(wire_switch_out_stage5[3]), .inData_4(wire_switch_out_stage5[4]), .inData_5(wire_switch_out_stage5[5]), .inData_6(wire_switch_out_stage5[6]), .inData_7(wire_switch_out_stage5[7]), .inData_8(wire_switch_out_stage5[8]), .inData_9(wire_switch_out_stage5[9]), .inData_10(wire_switch_out_stage5[10]), .inData_11(wire_switch_out_stage5[11]), .inData_12(wire_switch_out_stage5[12]), .inData_13(wire_switch_out_stage5[13]), .inData_14(wire_switch_out_stage5[14]), .inData_15(wire_switch_out_stage5[15]), .inData_16(wire_switch_out_stage5[16]), .inData_17(wire_switch_out_stage5[17]), .inData_18(wire_switch_out_stage5[18]), .inData_19(wire_switch_out_stage5[19]), .inData_20(wire_switch_out_stage5[20]), .inData_21(wire_switch_out_stage5[21]), .inData_22(wire_switch_out_stage5[22]), .inData_23(wire_switch_out_stage5[23]), .inData_24(wire_switch_out_stage5[24]), .inData_25(wire_switch_out_stage5[25]), .inData_26(wire_switch_out_stage5[26]), .inData_27(wire_switch_out_stage5[27]), .inData_28(wire_switch_out_stage5[28]), .inData_29(wire_switch_out_stage5[29]), .inData_30(wire_switch_out_stage5[30]), .inData_31(wire_switch_out_stage5[31]), .inData_32(wire_switch_out_stage5[32]), .inData_33(wire_switch_out_stage5[33]), .inData_34(wire_switch_out_stage5[34]), .inData_35(wire_switch_out_stage5[35]), .inData_36(wire_switch_out_stage5[36]), .inData_37(wire_switch_out_stage5[37]), .inData_38(wire_switch_out_stage5[38]), .inData_39(wire_switch_out_stage5[39]), .inData_40(wire_switch_out_stage5[40]), .inData_41(wire_switch_out_stage5[41]), .inData_42(wire_switch_out_stage5[42]), .inData_43(wire_switch_out_stage5[43]), .inData_44(wire_switch_out_stage5[44]), .inData_45(wire_switch_out_stage5[45]), .inData_46(wire_switch_out_stage5[46]), .inData_47(wire_switch_out_stage5[47]), .inData_48(wire_switch_out_stage5[48]), .inData_49(wire_switch_out_stage5[49]), .inData_50(wire_switch_out_stage5[50]), .inData_51(wire_switch_out_stage5[51]), .inData_52(wire_switch_out_stage5[52]), .inData_53(wire_switch_out_stage5[53]), .inData_54(wire_switch_out_stage5[54]), .inData_55(wire_switch_out_stage5[55]), .inData_56(wire_switch_out_stage5[56]), .inData_57(wire_switch_out_stage5[57]), .inData_58(wire_switch_out_stage5[58]), .inData_59(wire_switch_out_stage5[59]), .inData_60(wire_switch_out_stage5[60]), .inData_61(wire_switch_out_stage5[61]), .inData_62(wire_switch_out_stage5[62]), .inData_63(wire_switch_out_stage5[63]), .inData_64(wire_switch_out_stage5[64]), .inData_65(wire_switch_out_stage5[65]), .inData_66(wire_switch_out_stage5[66]), .inData_67(wire_switch_out_stage5[67]), .inData_68(wire_switch_out_stage5[68]), .inData_69(wire_switch_out_stage5[69]), .inData_70(wire_switch_out_stage5[70]), .inData_71(wire_switch_out_stage5[71]), .inData_72(wire_switch_out_stage5[72]), .inData_73(wire_switch_out_stage5[73]), .inData_74(wire_switch_out_stage5[74]), .inData_75(wire_switch_out_stage5[75]), .inData_76(wire_switch_out_stage5[76]), .inData_77(wire_switch_out_stage5[77]), .inData_78(wire_switch_out_stage5[78]), .inData_79(wire_switch_out_stage5[79]), .inData_80(wire_switch_out_stage5[80]), .inData_81(wire_switch_out_stage5[81]), .inData_82(wire_switch_out_stage5[82]), .inData_83(wire_switch_out_stage5[83]), .inData_84(wire_switch_out_stage5[84]), .inData_85(wire_switch_out_stage5[85]), .inData_86(wire_switch_out_stage5[86]), .inData_87(wire_switch_out_stage5[87]), .inData_88(wire_switch_out_stage5[88]), .inData_89(wire_switch_out_stage5[89]), .inData_90(wire_switch_out_stage5[90]), .inData_91(wire_switch_out_stage5[91]), .inData_92(wire_switch_out_stage5[92]), .inData_93(wire_switch_out_stage5[93]), .inData_94(wire_switch_out_stage5[94]), .inData_95(wire_switch_out_stage5[95]), .inData_96(wire_switch_out_stage5[96]), .inData_97(wire_switch_out_stage5[97]), .inData_98(wire_switch_out_stage5[98]), .inData_99(wire_switch_out_stage5[99]), .inData_100(wire_switch_out_stage5[100]), .inData_101(wire_switch_out_stage5[101]), .inData_102(wire_switch_out_stage5[102]), .inData_103(wire_switch_out_stage5[103]), .inData_104(wire_switch_out_stage5[104]), .inData_105(wire_switch_out_stage5[105]), .inData_106(wire_switch_out_stage5[106]), .inData_107(wire_switch_out_stage5[107]), .inData_108(wire_switch_out_stage5[108]), .inData_109(wire_switch_out_stage5[109]), .inData_110(wire_switch_out_stage5[110]), .inData_111(wire_switch_out_stage5[111]), .inData_112(wire_switch_out_stage5[112]), .inData_113(wire_switch_out_stage5[113]), .inData_114(wire_switch_out_stage5[114]), .inData_115(wire_switch_out_stage5[115]), .inData_116(wire_switch_out_stage5[116]), .inData_117(wire_switch_out_stage5[117]), .inData_118(wire_switch_out_stage5[118]), .inData_119(wire_switch_out_stage5[119]), .inData_120(wire_switch_out_stage5[120]), .inData_121(wire_switch_out_stage5[121]), .inData_122(wire_switch_out_stage5[122]), .inData_123(wire_switch_out_stage5[123]), .inData_124(wire_switch_out_stage5[124]), .inData_125(wire_switch_out_stage5[125]), .inData_126(wire_switch_out_stage5[126]), .inData_127(wire_switch_out_stage5[127]), .inData_128(wire_switch_out_stage5[128]), .inData_129(wire_switch_out_stage5[129]), .inData_130(wire_switch_out_stage5[130]), .inData_131(wire_switch_out_stage5[131]), .inData_132(wire_switch_out_stage5[132]), .inData_133(wire_switch_out_stage5[133]), .inData_134(wire_switch_out_stage5[134]), .inData_135(wire_switch_out_stage5[135]), .inData_136(wire_switch_out_stage5[136]), .inData_137(wire_switch_out_stage5[137]), .inData_138(wire_switch_out_stage5[138]), .inData_139(wire_switch_out_stage5[139]), .inData_140(wire_switch_out_stage5[140]), .inData_141(wire_switch_out_stage5[141]), .inData_142(wire_switch_out_stage5[142]), .inData_143(wire_switch_out_stage5[143]), .inData_144(wire_switch_out_stage5[144]), .inData_145(wire_switch_out_stage5[145]), .inData_146(wire_switch_out_stage5[146]), .inData_147(wire_switch_out_stage5[147]), .inData_148(wire_switch_out_stage5[148]), .inData_149(wire_switch_out_stage5[149]), .inData_150(wire_switch_out_stage5[150]), .inData_151(wire_switch_out_stage5[151]), .inData_152(wire_switch_out_stage5[152]), .inData_153(wire_switch_out_stage5[153]), .inData_154(wire_switch_out_stage5[154]), .inData_155(wire_switch_out_stage5[155]), .inData_156(wire_switch_out_stage5[156]), .inData_157(wire_switch_out_stage5[157]), .inData_158(wire_switch_out_stage5[158]), .inData_159(wire_switch_out_stage5[159]), .inData_160(wire_switch_out_stage5[160]), .inData_161(wire_switch_out_stage5[161]), .inData_162(wire_switch_out_stage5[162]), .inData_163(wire_switch_out_stage5[163]), .inData_164(wire_switch_out_stage5[164]), .inData_165(wire_switch_out_stage5[165]), .inData_166(wire_switch_out_stage5[166]), .inData_167(wire_switch_out_stage5[167]), .inData_168(wire_switch_out_stage5[168]), .inData_169(wire_switch_out_stage5[169]), .inData_170(wire_switch_out_stage5[170]), .inData_171(wire_switch_out_stage5[171]), .inData_172(wire_switch_out_stage5[172]), .inData_173(wire_switch_out_stage5[173]), .inData_174(wire_switch_out_stage5[174]), .inData_175(wire_switch_out_stage5[175]), .inData_176(wire_switch_out_stage5[176]), .inData_177(wire_switch_out_stage5[177]), .inData_178(wire_switch_out_stage5[178]), .inData_179(wire_switch_out_stage5[179]), .inData_180(wire_switch_out_stage5[180]), .inData_181(wire_switch_out_stage5[181]), .inData_182(wire_switch_out_stage5[182]), .inData_183(wire_switch_out_stage5[183]), .inData_184(wire_switch_out_stage5[184]), .inData_185(wire_switch_out_stage5[185]), .inData_186(wire_switch_out_stage5[186]), .inData_187(wire_switch_out_stage5[187]), .inData_188(wire_switch_out_stage5[188]), .inData_189(wire_switch_out_stage5[189]), .inData_190(wire_switch_out_stage5[190]), .inData_191(wire_switch_out_stage5[191]), .inData_192(wire_switch_out_stage5[192]), .inData_193(wire_switch_out_stage5[193]), .inData_194(wire_switch_out_stage5[194]), .inData_195(wire_switch_out_stage5[195]), .inData_196(wire_switch_out_stage5[196]), .inData_197(wire_switch_out_stage5[197]), .inData_198(wire_switch_out_stage5[198]), .inData_199(wire_switch_out_stage5[199]), .inData_200(wire_switch_out_stage5[200]), .inData_201(wire_switch_out_stage5[201]), .inData_202(wire_switch_out_stage5[202]), .inData_203(wire_switch_out_stage5[203]), .inData_204(wire_switch_out_stage5[204]), .inData_205(wire_switch_out_stage5[205]), .inData_206(wire_switch_out_stage5[206]), .inData_207(wire_switch_out_stage5[207]), .inData_208(wire_switch_out_stage5[208]), .inData_209(wire_switch_out_stage5[209]), .inData_210(wire_switch_out_stage5[210]), .inData_211(wire_switch_out_stage5[211]), .inData_212(wire_switch_out_stage5[212]), .inData_213(wire_switch_out_stage5[213]), .inData_214(wire_switch_out_stage5[214]), .inData_215(wire_switch_out_stage5[215]), .inData_216(wire_switch_out_stage5[216]), .inData_217(wire_switch_out_stage5[217]), .inData_218(wire_switch_out_stage5[218]), .inData_219(wire_switch_out_stage5[219]), .inData_220(wire_switch_out_stage5[220]), .inData_221(wire_switch_out_stage5[221]), .inData_222(wire_switch_out_stage5[222]), .inData_223(wire_switch_out_stage5[223]), .inData_224(wire_switch_out_stage5[224]), .inData_225(wire_switch_out_stage5[225]), .inData_226(wire_switch_out_stage5[226]), .inData_227(wire_switch_out_stage5[227]), .inData_228(wire_switch_out_stage5[228]), .inData_229(wire_switch_out_stage5[229]), .inData_230(wire_switch_out_stage5[230]), .inData_231(wire_switch_out_stage5[231]), .inData_232(wire_switch_out_stage5[232]), .inData_233(wire_switch_out_stage5[233]), .inData_234(wire_switch_out_stage5[234]), .inData_235(wire_switch_out_stage5[235]), .inData_236(wire_switch_out_stage5[236]), .inData_237(wire_switch_out_stage5[237]), .inData_238(wire_switch_out_stage5[238]), .inData_239(wire_switch_out_stage5[239]), .inData_240(wire_switch_out_stage5[240]), .inData_241(wire_switch_out_stage5[241]), .inData_242(wire_switch_out_stage5[242]), .inData_243(wire_switch_out_stage5[243]), .inData_244(wire_switch_out_stage5[244]), .inData_245(wire_switch_out_stage5[245]), .inData_246(wire_switch_out_stage5[246]), .inData_247(wire_switch_out_stage5[247]), .inData_248(wire_switch_out_stage5[248]), .inData_249(wire_switch_out_stage5[249]), .inData_250(wire_switch_out_stage5[250]), .inData_251(wire_switch_out_stage5[251]), .inData_252(wire_switch_out_stage5[252]), .inData_253(wire_switch_out_stage5[253]), .inData_254(wire_switch_out_stage5[254]), .inData_255(wire_switch_out_stage5[255]), 
        .outData_0(wire_switch_in_stage4[0]), .outData_1(wire_switch_in_stage4[1]), .outData_2(wire_switch_in_stage4[2]), .outData_3(wire_switch_in_stage4[3]), .outData_4(wire_switch_in_stage4[4]), .outData_5(wire_switch_in_stage4[5]), .outData_6(wire_switch_in_stage4[6]), .outData_7(wire_switch_in_stage4[7]), .outData_8(wire_switch_in_stage4[8]), .outData_9(wire_switch_in_stage4[9]), .outData_10(wire_switch_in_stage4[10]), .outData_11(wire_switch_in_stage4[11]), .outData_12(wire_switch_in_stage4[12]), .outData_13(wire_switch_in_stage4[13]), .outData_14(wire_switch_in_stage4[14]), .outData_15(wire_switch_in_stage4[15]), .outData_16(wire_switch_in_stage4[16]), .outData_17(wire_switch_in_stage4[17]), .outData_18(wire_switch_in_stage4[18]), .outData_19(wire_switch_in_stage4[19]), .outData_20(wire_switch_in_stage4[20]), .outData_21(wire_switch_in_stage4[21]), .outData_22(wire_switch_in_stage4[22]), .outData_23(wire_switch_in_stage4[23]), .outData_24(wire_switch_in_stage4[24]), .outData_25(wire_switch_in_stage4[25]), .outData_26(wire_switch_in_stage4[26]), .outData_27(wire_switch_in_stage4[27]), .outData_28(wire_switch_in_stage4[28]), .outData_29(wire_switch_in_stage4[29]), .outData_30(wire_switch_in_stage4[30]), .outData_31(wire_switch_in_stage4[31]), .outData_32(wire_switch_in_stage4[32]), .outData_33(wire_switch_in_stage4[33]), .outData_34(wire_switch_in_stage4[34]), .outData_35(wire_switch_in_stage4[35]), .outData_36(wire_switch_in_stage4[36]), .outData_37(wire_switch_in_stage4[37]), .outData_38(wire_switch_in_stage4[38]), .outData_39(wire_switch_in_stage4[39]), .outData_40(wire_switch_in_stage4[40]), .outData_41(wire_switch_in_stage4[41]), .outData_42(wire_switch_in_stage4[42]), .outData_43(wire_switch_in_stage4[43]), .outData_44(wire_switch_in_stage4[44]), .outData_45(wire_switch_in_stage4[45]), .outData_46(wire_switch_in_stage4[46]), .outData_47(wire_switch_in_stage4[47]), .outData_48(wire_switch_in_stage4[48]), .outData_49(wire_switch_in_stage4[49]), .outData_50(wire_switch_in_stage4[50]), .outData_51(wire_switch_in_stage4[51]), .outData_52(wire_switch_in_stage4[52]), .outData_53(wire_switch_in_stage4[53]), .outData_54(wire_switch_in_stage4[54]), .outData_55(wire_switch_in_stage4[55]), .outData_56(wire_switch_in_stage4[56]), .outData_57(wire_switch_in_stage4[57]), .outData_58(wire_switch_in_stage4[58]), .outData_59(wire_switch_in_stage4[59]), .outData_60(wire_switch_in_stage4[60]), .outData_61(wire_switch_in_stage4[61]), .outData_62(wire_switch_in_stage4[62]), .outData_63(wire_switch_in_stage4[63]), .outData_64(wire_switch_in_stage4[64]), .outData_65(wire_switch_in_stage4[65]), .outData_66(wire_switch_in_stage4[66]), .outData_67(wire_switch_in_stage4[67]), .outData_68(wire_switch_in_stage4[68]), .outData_69(wire_switch_in_stage4[69]), .outData_70(wire_switch_in_stage4[70]), .outData_71(wire_switch_in_stage4[71]), .outData_72(wire_switch_in_stage4[72]), .outData_73(wire_switch_in_stage4[73]), .outData_74(wire_switch_in_stage4[74]), .outData_75(wire_switch_in_stage4[75]), .outData_76(wire_switch_in_stage4[76]), .outData_77(wire_switch_in_stage4[77]), .outData_78(wire_switch_in_stage4[78]), .outData_79(wire_switch_in_stage4[79]), .outData_80(wire_switch_in_stage4[80]), .outData_81(wire_switch_in_stage4[81]), .outData_82(wire_switch_in_stage4[82]), .outData_83(wire_switch_in_stage4[83]), .outData_84(wire_switch_in_stage4[84]), .outData_85(wire_switch_in_stage4[85]), .outData_86(wire_switch_in_stage4[86]), .outData_87(wire_switch_in_stage4[87]), .outData_88(wire_switch_in_stage4[88]), .outData_89(wire_switch_in_stage4[89]), .outData_90(wire_switch_in_stage4[90]), .outData_91(wire_switch_in_stage4[91]), .outData_92(wire_switch_in_stage4[92]), .outData_93(wire_switch_in_stage4[93]), .outData_94(wire_switch_in_stage4[94]), .outData_95(wire_switch_in_stage4[95]), .outData_96(wire_switch_in_stage4[96]), .outData_97(wire_switch_in_stage4[97]), .outData_98(wire_switch_in_stage4[98]), .outData_99(wire_switch_in_stage4[99]), .outData_100(wire_switch_in_stage4[100]), .outData_101(wire_switch_in_stage4[101]), .outData_102(wire_switch_in_stage4[102]), .outData_103(wire_switch_in_stage4[103]), .outData_104(wire_switch_in_stage4[104]), .outData_105(wire_switch_in_stage4[105]), .outData_106(wire_switch_in_stage4[106]), .outData_107(wire_switch_in_stage4[107]), .outData_108(wire_switch_in_stage4[108]), .outData_109(wire_switch_in_stage4[109]), .outData_110(wire_switch_in_stage4[110]), .outData_111(wire_switch_in_stage4[111]), .outData_112(wire_switch_in_stage4[112]), .outData_113(wire_switch_in_stage4[113]), .outData_114(wire_switch_in_stage4[114]), .outData_115(wire_switch_in_stage4[115]), .outData_116(wire_switch_in_stage4[116]), .outData_117(wire_switch_in_stage4[117]), .outData_118(wire_switch_in_stage4[118]), .outData_119(wire_switch_in_stage4[119]), .outData_120(wire_switch_in_stage4[120]), .outData_121(wire_switch_in_stage4[121]), .outData_122(wire_switch_in_stage4[122]), .outData_123(wire_switch_in_stage4[123]), .outData_124(wire_switch_in_stage4[124]), .outData_125(wire_switch_in_stage4[125]), .outData_126(wire_switch_in_stage4[126]), .outData_127(wire_switch_in_stage4[127]), .outData_128(wire_switch_in_stage4[128]), .outData_129(wire_switch_in_stage4[129]), .outData_130(wire_switch_in_stage4[130]), .outData_131(wire_switch_in_stage4[131]), .outData_132(wire_switch_in_stage4[132]), .outData_133(wire_switch_in_stage4[133]), .outData_134(wire_switch_in_stage4[134]), .outData_135(wire_switch_in_stage4[135]), .outData_136(wire_switch_in_stage4[136]), .outData_137(wire_switch_in_stage4[137]), .outData_138(wire_switch_in_stage4[138]), .outData_139(wire_switch_in_stage4[139]), .outData_140(wire_switch_in_stage4[140]), .outData_141(wire_switch_in_stage4[141]), .outData_142(wire_switch_in_stage4[142]), .outData_143(wire_switch_in_stage4[143]), .outData_144(wire_switch_in_stage4[144]), .outData_145(wire_switch_in_stage4[145]), .outData_146(wire_switch_in_stage4[146]), .outData_147(wire_switch_in_stage4[147]), .outData_148(wire_switch_in_stage4[148]), .outData_149(wire_switch_in_stage4[149]), .outData_150(wire_switch_in_stage4[150]), .outData_151(wire_switch_in_stage4[151]), .outData_152(wire_switch_in_stage4[152]), .outData_153(wire_switch_in_stage4[153]), .outData_154(wire_switch_in_stage4[154]), .outData_155(wire_switch_in_stage4[155]), .outData_156(wire_switch_in_stage4[156]), .outData_157(wire_switch_in_stage4[157]), .outData_158(wire_switch_in_stage4[158]), .outData_159(wire_switch_in_stage4[159]), .outData_160(wire_switch_in_stage4[160]), .outData_161(wire_switch_in_stage4[161]), .outData_162(wire_switch_in_stage4[162]), .outData_163(wire_switch_in_stage4[163]), .outData_164(wire_switch_in_stage4[164]), .outData_165(wire_switch_in_stage4[165]), .outData_166(wire_switch_in_stage4[166]), .outData_167(wire_switch_in_stage4[167]), .outData_168(wire_switch_in_stage4[168]), .outData_169(wire_switch_in_stage4[169]), .outData_170(wire_switch_in_stage4[170]), .outData_171(wire_switch_in_stage4[171]), .outData_172(wire_switch_in_stage4[172]), .outData_173(wire_switch_in_stage4[173]), .outData_174(wire_switch_in_stage4[174]), .outData_175(wire_switch_in_stage4[175]), .outData_176(wire_switch_in_stage4[176]), .outData_177(wire_switch_in_stage4[177]), .outData_178(wire_switch_in_stage4[178]), .outData_179(wire_switch_in_stage4[179]), .outData_180(wire_switch_in_stage4[180]), .outData_181(wire_switch_in_stage4[181]), .outData_182(wire_switch_in_stage4[182]), .outData_183(wire_switch_in_stage4[183]), .outData_184(wire_switch_in_stage4[184]), .outData_185(wire_switch_in_stage4[185]), .outData_186(wire_switch_in_stage4[186]), .outData_187(wire_switch_in_stage4[187]), .outData_188(wire_switch_in_stage4[188]), .outData_189(wire_switch_in_stage4[189]), .outData_190(wire_switch_in_stage4[190]), .outData_191(wire_switch_in_stage4[191]), .outData_192(wire_switch_in_stage4[192]), .outData_193(wire_switch_in_stage4[193]), .outData_194(wire_switch_in_stage4[194]), .outData_195(wire_switch_in_stage4[195]), .outData_196(wire_switch_in_stage4[196]), .outData_197(wire_switch_in_stage4[197]), .outData_198(wire_switch_in_stage4[198]), .outData_199(wire_switch_in_stage4[199]), .outData_200(wire_switch_in_stage4[200]), .outData_201(wire_switch_in_stage4[201]), .outData_202(wire_switch_in_stage4[202]), .outData_203(wire_switch_in_stage4[203]), .outData_204(wire_switch_in_stage4[204]), .outData_205(wire_switch_in_stage4[205]), .outData_206(wire_switch_in_stage4[206]), .outData_207(wire_switch_in_stage4[207]), .outData_208(wire_switch_in_stage4[208]), .outData_209(wire_switch_in_stage4[209]), .outData_210(wire_switch_in_stage4[210]), .outData_211(wire_switch_in_stage4[211]), .outData_212(wire_switch_in_stage4[212]), .outData_213(wire_switch_in_stage4[213]), .outData_214(wire_switch_in_stage4[214]), .outData_215(wire_switch_in_stage4[215]), .outData_216(wire_switch_in_stage4[216]), .outData_217(wire_switch_in_stage4[217]), .outData_218(wire_switch_in_stage4[218]), .outData_219(wire_switch_in_stage4[219]), .outData_220(wire_switch_in_stage4[220]), .outData_221(wire_switch_in_stage4[221]), .outData_222(wire_switch_in_stage4[222]), .outData_223(wire_switch_in_stage4[223]), .outData_224(wire_switch_in_stage4[224]), .outData_225(wire_switch_in_stage4[225]), .outData_226(wire_switch_in_stage4[226]), .outData_227(wire_switch_in_stage4[227]), .outData_228(wire_switch_in_stage4[228]), .outData_229(wire_switch_in_stage4[229]), .outData_230(wire_switch_in_stage4[230]), .outData_231(wire_switch_in_stage4[231]), .outData_232(wire_switch_in_stage4[232]), .outData_233(wire_switch_in_stage4[233]), .outData_234(wire_switch_in_stage4[234]), .outData_235(wire_switch_in_stage4[235]), .outData_236(wire_switch_in_stage4[236]), .outData_237(wire_switch_in_stage4[237]), .outData_238(wire_switch_in_stage4[238]), .outData_239(wire_switch_in_stage4[239]), .outData_240(wire_switch_in_stage4[240]), .outData_241(wire_switch_in_stage4[241]), .outData_242(wire_switch_in_stage4[242]), .outData_243(wire_switch_in_stage4[243]), .outData_244(wire_switch_in_stage4[244]), .outData_245(wire_switch_in_stage4[245]), .outData_246(wire_switch_in_stage4[246]), .outData_247(wire_switch_in_stage4[247]), .outData_248(wire_switch_in_stage4[248]), .outData_249(wire_switch_in_stage4[249]), .outData_250(wire_switch_in_stage4[250]), .outData_251(wire_switch_in_stage4[251]), .outData_252(wire_switch_in_stage4[252]), .outData_253(wire_switch_in_stage4[253]), .outData_254(wire_switch_in_stage4[254]), .outData_255(wire_switch_in_stage4[255]), 
        .in_start(in_start_stage4), .out_start(con_in_start_stage4), .clk(clk), .rst(rst)); 

  
  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[0] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[1] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[2] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[3] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[4] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[5] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[6] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[7] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[8] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[9] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[10] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[11] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[12] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[13] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[14] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[15] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[16] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[17] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[18] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[19] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[20] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[21] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[22] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[23] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[24] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[25] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[26] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[27] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[28] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[29] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[30] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[31] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[32] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[33] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[34] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[35] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[36] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[37] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[38] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[39] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[40] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[41] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[42] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[43] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[44] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[45] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[46] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[47] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[48] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[49] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[50] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[51] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[52] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[53] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[54] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[55] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[56] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[57] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[58] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[59] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[60] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[61] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[62] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[63] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[64] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[65] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[66] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[67] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[68] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[69] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[70] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[71] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[72] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[73] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[74] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[75] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[76] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[77] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[78] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[79] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[80] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[81] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[82] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[83] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[84] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[85] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[86] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[87] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[88] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[89] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[90] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[91] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[92] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[93] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[94] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[95] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[96] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[97] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[98] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[99] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[100] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[101] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[102] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[103] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[104] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[105] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[106] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[107] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[108] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[109] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[110] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[111] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[112] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[113] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[114] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[115] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[116] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[117] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[118] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[119] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[120] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[121] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[122] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[123] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[124] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[125] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[126] <= counter_w[3]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage4[127] <= counter_w[3]; 
  end                            

  wire [DATA_WIDTH-1:0] wire_switch_in_stage3[255:0];
  wire [DATA_WIDTH-1:0] wire_switch_out_stage3[255:0];
  reg [127:0] wire_ctrl_stage3;

  switches_stage_st3_0_R switch_stage_3(
        .inData_0(wire_switch_in_stage3[0]), .inData_1(wire_switch_in_stage3[1]), .inData_2(wire_switch_in_stage3[2]), .inData_3(wire_switch_in_stage3[3]), .inData_4(wire_switch_in_stage3[4]), .inData_5(wire_switch_in_stage3[5]), .inData_6(wire_switch_in_stage3[6]), .inData_7(wire_switch_in_stage3[7]), .inData_8(wire_switch_in_stage3[8]), .inData_9(wire_switch_in_stage3[9]), .inData_10(wire_switch_in_stage3[10]), .inData_11(wire_switch_in_stage3[11]), .inData_12(wire_switch_in_stage3[12]), .inData_13(wire_switch_in_stage3[13]), .inData_14(wire_switch_in_stage3[14]), .inData_15(wire_switch_in_stage3[15]), .inData_16(wire_switch_in_stage3[16]), .inData_17(wire_switch_in_stage3[17]), .inData_18(wire_switch_in_stage3[18]), .inData_19(wire_switch_in_stage3[19]), .inData_20(wire_switch_in_stage3[20]), .inData_21(wire_switch_in_stage3[21]), .inData_22(wire_switch_in_stage3[22]), .inData_23(wire_switch_in_stage3[23]), .inData_24(wire_switch_in_stage3[24]), .inData_25(wire_switch_in_stage3[25]), .inData_26(wire_switch_in_stage3[26]), .inData_27(wire_switch_in_stage3[27]), .inData_28(wire_switch_in_stage3[28]), .inData_29(wire_switch_in_stage3[29]), .inData_30(wire_switch_in_stage3[30]), .inData_31(wire_switch_in_stage3[31]), .inData_32(wire_switch_in_stage3[32]), .inData_33(wire_switch_in_stage3[33]), .inData_34(wire_switch_in_stage3[34]), .inData_35(wire_switch_in_stage3[35]), .inData_36(wire_switch_in_stage3[36]), .inData_37(wire_switch_in_stage3[37]), .inData_38(wire_switch_in_stage3[38]), .inData_39(wire_switch_in_stage3[39]), .inData_40(wire_switch_in_stage3[40]), .inData_41(wire_switch_in_stage3[41]), .inData_42(wire_switch_in_stage3[42]), .inData_43(wire_switch_in_stage3[43]), .inData_44(wire_switch_in_stage3[44]), .inData_45(wire_switch_in_stage3[45]), .inData_46(wire_switch_in_stage3[46]), .inData_47(wire_switch_in_stage3[47]), .inData_48(wire_switch_in_stage3[48]), .inData_49(wire_switch_in_stage3[49]), .inData_50(wire_switch_in_stage3[50]), .inData_51(wire_switch_in_stage3[51]), .inData_52(wire_switch_in_stage3[52]), .inData_53(wire_switch_in_stage3[53]), .inData_54(wire_switch_in_stage3[54]), .inData_55(wire_switch_in_stage3[55]), .inData_56(wire_switch_in_stage3[56]), .inData_57(wire_switch_in_stage3[57]), .inData_58(wire_switch_in_stage3[58]), .inData_59(wire_switch_in_stage3[59]), .inData_60(wire_switch_in_stage3[60]), .inData_61(wire_switch_in_stage3[61]), .inData_62(wire_switch_in_stage3[62]), .inData_63(wire_switch_in_stage3[63]), .inData_64(wire_switch_in_stage3[64]), .inData_65(wire_switch_in_stage3[65]), .inData_66(wire_switch_in_stage3[66]), .inData_67(wire_switch_in_stage3[67]), .inData_68(wire_switch_in_stage3[68]), .inData_69(wire_switch_in_stage3[69]), .inData_70(wire_switch_in_stage3[70]), .inData_71(wire_switch_in_stage3[71]), .inData_72(wire_switch_in_stage3[72]), .inData_73(wire_switch_in_stage3[73]), .inData_74(wire_switch_in_stage3[74]), .inData_75(wire_switch_in_stage3[75]), .inData_76(wire_switch_in_stage3[76]), .inData_77(wire_switch_in_stage3[77]), .inData_78(wire_switch_in_stage3[78]), .inData_79(wire_switch_in_stage3[79]), .inData_80(wire_switch_in_stage3[80]), .inData_81(wire_switch_in_stage3[81]), .inData_82(wire_switch_in_stage3[82]), .inData_83(wire_switch_in_stage3[83]), .inData_84(wire_switch_in_stage3[84]), .inData_85(wire_switch_in_stage3[85]), .inData_86(wire_switch_in_stage3[86]), .inData_87(wire_switch_in_stage3[87]), .inData_88(wire_switch_in_stage3[88]), .inData_89(wire_switch_in_stage3[89]), .inData_90(wire_switch_in_stage3[90]), .inData_91(wire_switch_in_stage3[91]), .inData_92(wire_switch_in_stage3[92]), .inData_93(wire_switch_in_stage3[93]), .inData_94(wire_switch_in_stage3[94]), .inData_95(wire_switch_in_stage3[95]), .inData_96(wire_switch_in_stage3[96]), .inData_97(wire_switch_in_stage3[97]), .inData_98(wire_switch_in_stage3[98]), .inData_99(wire_switch_in_stage3[99]), .inData_100(wire_switch_in_stage3[100]), .inData_101(wire_switch_in_stage3[101]), .inData_102(wire_switch_in_stage3[102]), .inData_103(wire_switch_in_stage3[103]), .inData_104(wire_switch_in_stage3[104]), .inData_105(wire_switch_in_stage3[105]), .inData_106(wire_switch_in_stage3[106]), .inData_107(wire_switch_in_stage3[107]), .inData_108(wire_switch_in_stage3[108]), .inData_109(wire_switch_in_stage3[109]), .inData_110(wire_switch_in_stage3[110]), .inData_111(wire_switch_in_stage3[111]), .inData_112(wire_switch_in_stage3[112]), .inData_113(wire_switch_in_stage3[113]), .inData_114(wire_switch_in_stage3[114]), .inData_115(wire_switch_in_stage3[115]), .inData_116(wire_switch_in_stage3[116]), .inData_117(wire_switch_in_stage3[117]), .inData_118(wire_switch_in_stage3[118]), .inData_119(wire_switch_in_stage3[119]), .inData_120(wire_switch_in_stage3[120]), .inData_121(wire_switch_in_stage3[121]), .inData_122(wire_switch_in_stage3[122]), .inData_123(wire_switch_in_stage3[123]), .inData_124(wire_switch_in_stage3[124]), .inData_125(wire_switch_in_stage3[125]), .inData_126(wire_switch_in_stage3[126]), .inData_127(wire_switch_in_stage3[127]), .inData_128(wire_switch_in_stage3[128]), .inData_129(wire_switch_in_stage3[129]), .inData_130(wire_switch_in_stage3[130]), .inData_131(wire_switch_in_stage3[131]), .inData_132(wire_switch_in_stage3[132]), .inData_133(wire_switch_in_stage3[133]), .inData_134(wire_switch_in_stage3[134]), .inData_135(wire_switch_in_stage3[135]), .inData_136(wire_switch_in_stage3[136]), .inData_137(wire_switch_in_stage3[137]), .inData_138(wire_switch_in_stage3[138]), .inData_139(wire_switch_in_stage3[139]), .inData_140(wire_switch_in_stage3[140]), .inData_141(wire_switch_in_stage3[141]), .inData_142(wire_switch_in_stage3[142]), .inData_143(wire_switch_in_stage3[143]), .inData_144(wire_switch_in_stage3[144]), .inData_145(wire_switch_in_stage3[145]), .inData_146(wire_switch_in_stage3[146]), .inData_147(wire_switch_in_stage3[147]), .inData_148(wire_switch_in_stage3[148]), .inData_149(wire_switch_in_stage3[149]), .inData_150(wire_switch_in_stage3[150]), .inData_151(wire_switch_in_stage3[151]), .inData_152(wire_switch_in_stage3[152]), .inData_153(wire_switch_in_stage3[153]), .inData_154(wire_switch_in_stage3[154]), .inData_155(wire_switch_in_stage3[155]), .inData_156(wire_switch_in_stage3[156]), .inData_157(wire_switch_in_stage3[157]), .inData_158(wire_switch_in_stage3[158]), .inData_159(wire_switch_in_stage3[159]), .inData_160(wire_switch_in_stage3[160]), .inData_161(wire_switch_in_stage3[161]), .inData_162(wire_switch_in_stage3[162]), .inData_163(wire_switch_in_stage3[163]), .inData_164(wire_switch_in_stage3[164]), .inData_165(wire_switch_in_stage3[165]), .inData_166(wire_switch_in_stage3[166]), .inData_167(wire_switch_in_stage3[167]), .inData_168(wire_switch_in_stage3[168]), .inData_169(wire_switch_in_stage3[169]), .inData_170(wire_switch_in_stage3[170]), .inData_171(wire_switch_in_stage3[171]), .inData_172(wire_switch_in_stage3[172]), .inData_173(wire_switch_in_stage3[173]), .inData_174(wire_switch_in_stage3[174]), .inData_175(wire_switch_in_stage3[175]), .inData_176(wire_switch_in_stage3[176]), .inData_177(wire_switch_in_stage3[177]), .inData_178(wire_switch_in_stage3[178]), .inData_179(wire_switch_in_stage3[179]), .inData_180(wire_switch_in_stage3[180]), .inData_181(wire_switch_in_stage3[181]), .inData_182(wire_switch_in_stage3[182]), .inData_183(wire_switch_in_stage3[183]), .inData_184(wire_switch_in_stage3[184]), .inData_185(wire_switch_in_stage3[185]), .inData_186(wire_switch_in_stage3[186]), .inData_187(wire_switch_in_stage3[187]), .inData_188(wire_switch_in_stage3[188]), .inData_189(wire_switch_in_stage3[189]), .inData_190(wire_switch_in_stage3[190]), .inData_191(wire_switch_in_stage3[191]), .inData_192(wire_switch_in_stage3[192]), .inData_193(wire_switch_in_stage3[193]), .inData_194(wire_switch_in_stage3[194]), .inData_195(wire_switch_in_stage3[195]), .inData_196(wire_switch_in_stage3[196]), .inData_197(wire_switch_in_stage3[197]), .inData_198(wire_switch_in_stage3[198]), .inData_199(wire_switch_in_stage3[199]), .inData_200(wire_switch_in_stage3[200]), .inData_201(wire_switch_in_stage3[201]), .inData_202(wire_switch_in_stage3[202]), .inData_203(wire_switch_in_stage3[203]), .inData_204(wire_switch_in_stage3[204]), .inData_205(wire_switch_in_stage3[205]), .inData_206(wire_switch_in_stage3[206]), .inData_207(wire_switch_in_stage3[207]), .inData_208(wire_switch_in_stage3[208]), .inData_209(wire_switch_in_stage3[209]), .inData_210(wire_switch_in_stage3[210]), .inData_211(wire_switch_in_stage3[211]), .inData_212(wire_switch_in_stage3[212]), .inData_213(wire_switch_in_stage3[213]), .inData_214(wire_switch_in_stage3[214]), .inData_215(wire_switch_in_stage3[215]), .inData_216(wire_switch_in_stage3[216]), .inData_217(wire_switch_in_stage3[217]), .inData_218(wire_switch_in_stage3[218]), .inData_219(wire_switch_in_stage3[219]), .inData_220(wire_switch_in_stage3[220]), .inData_221(wire_switch_in_stage3[221]), .inData_222(wire_switch_in_stage3[222]), .inData_223(wire_switch_in_stage3[223]), .inData_224(wire_switch_in_stage3[224]), .inData_225(wire_switch_in_stage3[225]), .inData_226(wire_switch_in_stage3[226]), .inData_227(wire_switch_in_stage3[227]), .inData_228(wire_switch_in_stage3[228]), .inData_229(wire_switch_in_stage3[229]), .inData_230(wire_switch_in_stage3[230]), .inData_231(wire_switch_in_stage3[231]), .inData_232(wire_switch_in_stage3[232]), .inData_233(wire_switch_in_stage3[233]), .inData_234(wire_switch_in_stage3[234]), .inData_235(wire_switch_in_stage3[235]), .inData_236(wire_switch_in_stage3[236]), .inData_237(wire_switch_in_stage3[237]), .inData_238(wire_switch_in_stage3[238]), .inData_239(wire_switch_in_stage3[239]), .inData_240(wire_switch_in_stage3[240]), .inData_241(wire_switch_in_stage3[241]), .inData_242(wire_switch_in_stage3[242]), .inData_243(wire_switch_in_stage3[243]), .inData_244(wire_switch_in_stage3[244]), .inData_245(wire_switch_in_stage3[245]), .inData_246(wire_switch_in_stage3[246]), .inData_247(wire_switch_in_stage3[247]), .inData_248(wire_switch_in_stage3[248]), .inData_249(wire_switch_in_stage3[249]), .inData_250(wire_switch_in_stage3[250]), .inData_251(wire_switch_in_stage3[251]), .inData_252(wire_switch_in_stage3[252]), .inData_253(wire_switch_in_stage3[253]), .inData_254(wire_switch_in_stage3[254]), .inData_255(wire_switch_in_stage3[255]), 
        .outData_0(wire_switch_out_stage3[0]), .outData_1(wire_switch_out_stage3[1]), .outData_2(wire_switch_out_stage3[2]), .outData_3(wire_switch_out_stage3[3]), .outData_4(wire_switch_out_stage3[4]), .outData_5(wire_switch_out_stage3[5]), .outData_6(wire_switch_out_stage3[6]), .outData_7(wire_switch_out_stage3[7]), .outData_8(wire_switch_out_stage3[8]), .outData_9(wire_switch_out_stage3[9]), .outData_10(wire_switch_out_stage3[10]), .outData_11(wire_switch_out_stage3[11]), .outData_12(wire_switch_out_stage3[12]), .outData_13(wire_switch_out_stage3[13]), .outData_14(wire_switch_out_stage3[14]), .outData_15(wire_switch_out_stage3[15]), .outData_16(wire_switch_out_stage3[16]), .outData_17(wire_switch_out_stage3[17]), .outData_18(wire_switch_out_stage3[18]), .outData_19(wire_switch_out_stage3[19]), .outData_20(wire_switch_out_stage3[20]), .outData_21(wire_switch_out_stage3[21]), .outData_22(wire_switch_out_stage3[22]), .outData_23(wire_switch_out_stage3[23]), .outData_24(wire_switch_out_stage3[24]), .outData_25(wire_switch_out_stage3[25]), .outData_26(wire_switch_out_stage3[26]), .outData_27(wire_switch_out_stage3[27]), .outData_28(wire_switch_out_stage3[28]), .outData_29(wire_switch_out_stage3[29]), .outData_30(wire_switch_out_stage3[30]), .outData_31(wire_switch_out_stage3[31]), .outData_32(wire_switch_out_stage3[32]), .outData_33(wire_switch_out_stage3[33]), .outData_34(wire_switch_out_stage3[34]), .outData_35(wire_switch_out_stage3[35]), .outData_36(wire_switch_out_stage3[36]), .outData_37(wire_switch_out_stage3[37]), .outData_38(wire_switch_out_stage3[38]), .outData_39(wire_switch_out_stage3[39]), .outData_40(wire_switch_out_stage3[40]), .outData_41(wire_switch_out_stage3[41]), .outData_42(wire_switch_out_stage3[42]), .outData_43(wire_switch_out_stage3[43]), .outData_44(wire_switch_out_stage3[44]), .outData_45(wire_switch_out_stage3[45]), .outData_46(wire_switch_out_stage3[46]), .outData_47(wire_switch_out_stage3[47]), .outData_48(wire_switch_out_stage3[48]), .outData_49(wire_switch_out_stage3[49]), .outData_50(wire_switch_out_stage3[50]), .outData_51(wire_switch_out_stage3[51]), .outData_52(wire_switch_out_stage3[52]), .outData_53(wire_switch_out_stage3[53]), .outData_54(wire_switch_out_stage3[54]), .outData_55(wire_switch_out_stage3[55]), .outData_56(wire_switch_out_stage3[56]), .outData_57(wire_switch_out_stage3[57]), .outData_58(wire_switch_out_stage3[58]), .outData_59(wire_switch_out_stage3[59]), .outData_60(wire_switch_out_stage3[60]), .outData_61(wire_switch_out_stage3[61]), .outData_62(wire_switch_out_stage3[62]), .outData_63(wire_switch_out_stage3[63]), .outData_64(wire_switch_out_stage3[64]), .outData_65(wire_switch_out_stage3[65]), .outData_66(wire_switch_out_stage3[66]), .outData_67(wire_switch_out_stage3[67]), .outData_68(wire_switch_out_stage3[68]), .outData_69(wire_switch_out_stage3[69]), .outData_70(wire_switch_out_stage3[70]), .outData_71(wire_switch_out_stage3[71]), .outData_72(wire_switch_out_stage3[72]), .outData_73(wire_switch_out_stage3[73]), .outData_74(wire_switch_out_stage3[74]), .outData_75(wire_switch_out_stage3[75]), .outData_76(wire_switch_out_stage3[76]), .outData_77(wire_switch_out_stage3[77]), .outData_78(wire_switch_out_stage3[78]), .outData_79(wire_switch_out_stage3[79]), .outData_80(wire_switch_out_stage3[80]), .outData_81(wire_switch_out_stage3[81]), .outData_82(wire_switch_out_stage3[82]), .outData_83(wire_switch_out_stage3[83]), .outData_84(wire_switch_out_stage3[84]), .outData_85(wire_switch_out_stage3[85]), .outData_86(wire_switch_out_stage3[86]), .outData_87(wire_switch_out_stage3[87]), .outData_88(wire_switch_out_stage3[88]), .outData_89(wire_switch_out_stage3[89]), .outData_90(wire_switch_out_stage3[90]), .outData_91(wire_switch_out_stage3[91]), .outData_92(wire_switch_out_stage3[92]), .outData_93(wire_switch_out_stage3[93]), .outData_94(wire_switch_out_stage3[94]), .outData_95(wire_switch_out_stage3[95]), .outData_96(wire_switch_out_stage3[96]), .outData_97(wire_switch_out_stage3[97]), .outData_98(wire_switch_out_stage3[98]), .outData_99(wire_switch_out_stage3[99]), .outData_100(wire_switch_out_stage3[100]), .outData_101(wire_switch_out_stage3[101]), .outData_102(wire_switch_out_stage3[102]), .outData_103(wire_switch_out_stage3[103]), .outData_104(wire_switch_out_stage3[104]), .outData_105(wire_switch_out_stage3[105]), .outData_106(wire_switch_out_stage3[106]), .outData_107(wire_switch_out_stage3[107]), .outData_108(wire_switch_out_stage3[108]), .outData_109(wire_switch_out_stage3[109]), .outData_110(wire_switch_out_stage3[110]), .outData_111(wire_switch_out_stage3[111]), .outData_112(wire_switch_out_stage3[112]), .outData_113(wire_switch_out_stage3[113]), .outData_114(wire_switch_out_stage3[114]), .outData_115(wire_switch_out_stage3[115]), .outData_116(wire_switch_out_stage3[116]), .outData_117(wire_switch_out_stage3[117]), .outData_118(wire_switch_out_stage3[118]), .outData_119(wire_switch_out_stage3[119]), .outData_120(wire_switch_out_stage3[120]), .outData_121(wire_switch_out_stage3[121]), .outData_122(wire_switch_out_stage3[122]), .outData_123(wire_switch_out_stage3[123]), .outData_124(wire_switch_out_stage3[124]), .outData_125(wire_switch_out_stage3[125]), .outData_126(wire_switch_out_stage3[126]), .outData_127(wire_switch_out_stage3[127]), .outData_128(wire_switch_out_stage3[128]), .outData_129(wire_switch_out_stage3[129]), .outData_130(wire_switch_out_stage3[130]), .outData_131(wire_switch_out_stage3[131]), .outData_132(wire_switch_out_stage3[132]), .outData_133(wire_switch_out_stage3[133]), .outData_134(wire_switch_out_stage3[134]), .outData_135(wire_switch_out_stage3[135]), .outData_136(wire_switch_out_stage3[136]), .outData_137(wire_switch_out_stage3[137]), .outData_138(wire_switch_out_stage3[138]), .outData_139(wire_switch_out_stage3[139]), .outData_140(wire_switch_out_stage3[140]), .outData_141(wire_switch_out_stage3[141]), .outData_142(wire_switch_out_stage3[142]), .outData_143(wire_switch_out_stage3[143]), .outData_144(wire_switch_out_stage3[144]), .outData_145(wire_switch_out_stage3[145]), .outData_146(wire_switch_out_stage3[146]), .outData_147(wire_switch_out_stage3[147]), .outData_148(wire_switch_out_stage3[148]), .outData_149(wire_switch_out_stage3[149]), .outData_150(wire_switch_out_stage3[150]), .outData_151(wire_switch_out_stage3[151]), .outData_152(wire_switch_out_stage3[152]), .outData_153(wire_switch_out_stage3[153]), .outData_154(wire_switch_out_stage3[154]), .outData_155(wire_switch_out_stage3[155]), .outData_156(wire_switch_out_stage3[156]), .outData_157(wire_switch_out_stage3[157]), .outData_158(wire_switch_out_stage3[158]), .outData_159(wire_switch_out_stage3[159]), .outData_160(wire_switch_out_stage3[160]), .outData_161(wire_switch_out_stage3[161]), .outData_162(wire_switch_out_stage3[162]), .outData_163(wire_switch_out_stage3[163]), .outData_164(wire_switch_out_stage3[164]), .outData_165(wire_switch_out_stage3[165]), .outData_166(wire_switch_out_stage3[166]), .outData_167(wire_switch_out_stage3[167]), .outData_168(wire_switch_out_stage3[168]), .outData_169(wire_switch_out_stage3[169]), .outData_170(wire_switch_out_stage3[170]), .outData_171(wire_switch_out_stage3[171]), .outData_172(wire_switch_out_stage3[172]), .outData_173(wire_switch_out_stage3[173]), .outData_174(wire_switch_out_stage3[174]), .outData_175(wire_switch_out_stage3[175]), .outData_176(wire_switch_out_stage3[176]), .outData_177(wire_switch_out_stage3[177]), .outData_178(wire_switch_out_stage3[178]), .outData_179(wire_switch_out_stage3[179]), .outData_180(wire_switch_out_stage3[180]), .outData_181(wire_switch_out_stage3[181]), .outData_182(wire_switch_out_stage3[182]), .outData_183(wire_switch_out_stage3[183]), .outData_184(wire_switch_out_stage3[184]), .outData_185(wire_switch_out_stage3[185]), .outData_186(wire_switch_out_stage3[186]), .outData_187(wire_switch_out_stage3[187]), .outData_188(wire_switch_out_stage3[188]), .outData_189(wire_switch_out_stage3[189]), .outData_190(wire_switch_out_stage3[190]), .outData_191(wire_switch_out_stage3[191]), .outData_192(wire_switch_out_stage3[192]), .outData_193(wire_switch_out_stage3[193]), .outData_194(wire_switch_out_stage3[194]), .outData_195(wire_switch_out_stage3[195]), .outData_196(wire_switch_out_stage3[196]), .outData_197(wire_switch_out_stage3[197]), .outData_198(wire_switch_out_stage3[198]), .outData_199(wire_switch_out_stage3[199]), .outData_200(wire_switch_out_stage3[200]), .outData_201(wire_switch_out_stage3[201]), .outData_202(wire_switch_out_stage3[202]), .outData_203(wire_switch_out_stage3[203]), .outData_204(wire_switch_out_stage3[204]), .outData_205(wire_switch_out_stage3[205]), .outData_206(wire_switch_out_stage3[206]), .outData_207(wire_switch_out_stage3[207]), .outData_208(wire_switch_out_stage3[208]), .outData_209(wire_switch_out_stage3[209]), .outData_210(wire_switch_out_stage3[210]), .outData_211(wire_switch_out_stage3[211]), .outData_212(wire_switch_out_stage3[212]), .outData_213(wire_switch_out_stage3[213]), .outData_214(wire_switch_out_stage3[214]), .outData_215(wire_switch_out_stage3[215]), .outData_216(wire_switch_out_stage3[216]), .outData_217(wire_switch_out_stage3[217]), .outData_218(wire_switch_out_stage3[218]), .outData_219(wire_switch_out_stage3[219]), .outData_220(wire_switch_out_stage3[220]), .outData_221(wire_switch_out_stage3[221]), .outData_222(wire_switch_out_stage3[222]), .outData_223(wire_switch_out_stage3[223]), .outData_224(wire_switch_out_stage3[224]), .outData_225(wire_switch_out_stage3[225]), .outData_226(wire_switch_out_stage3[226]), .outData_227(wire_switch_out_stage3[227]), .outData_228(wire_switch_out_stage3[228]), .outData_229(wire_switch_out_stage3[229]), .outData_230(wire_switch_out_stage3[230]), .outData_231(wire_switch_out_stage3[231]), .outData_232(wire_switch_out_stage3[232]), .outData_233(wire_switch_out_stage3[233]), .outData_234(wire_switch_out_stage3[234]), .outData_235(wire_switch_out_stage3[235]), .outData_236(wire_switch_out_stage3[236]), .outData_237(wire_switch_out_stage3[237]), .outData_238(wire_switch_out_stage3[238]), .outData_239(wire_switch_out_stage3[239]), .outData_240(wire_switch_out_stage3[240]), .outData_241(wire_switch_out_stage3[241]), .outData_242(wire_switch_out_stage3[242]), .outData_243(wire_switch_out_stage3[243]), .outData_244(wire_switch_out_stage3[244]), .outData_245(wire_switch_out_stage3[245]), .outData_246(wire_switch_out_stage3[246]), .outData_247(wire_switch_out_stage3[247]), .outData_248(wire_switch_out_stage3[248]), .outData_249(wire_switch_out_stage3[249]), .outData_250(wire_switch_out_stage3[250]), .outData_251(wire_switch_out_stage3[251]), .outData_252(wire_switch_out_stage3[252]), .outData_253(wire_switch_out_stage3[253]), .outData_254(wire_switch_out_stage3[254]), .outData_255(wire_switch_out_stage3[255]), 
        .in_start(con_in_start_stage3), .out_start(in_start_stage2), .ctrl(wire_ctrl_stage3), .clk(clk), .rst(rst));
  
  wireCon_dp256_st3_R wire_stage_3(
        .inData_0(wire_switch_out_stage4[0]), .inData_1(wire_switch_out_stage4[1]), .inData_2(wire_switch_out_stage4[2]), .inData_3(wire_switch_out_stage4[3]), .inData_4(wire_switch_out_stage4[4]), .inData_5(wire_switch_out_stage4[5]), .inData_6(wire_switch_out_stage4[6]), .inData_7(wire_switch_out_stage4[7]), .inData_8(wire_switch_out_stage4[8]), .inData_9(wire_switch_out_stage4[9]), .inData_10(wire_switch_out_stage4[10]), .inData_11(wire_switch_out_stage4[11]), .inData_12(wire_switch_out_stage4[12]), .inData_13(wire_switch_out_stage4[13]), .inData_14(wire_switch_out_stage4[14]), .inData_15(wire_switch_out_stage4[15]), .inData_16(wire_switch_out_stage4[16]), .inData_17(wire_switch_out_stage4[17]), .inData_18(wire_switch_out_stage4[18]), .inData_19(wire_switch_out_stage4[19]), .inData_20(wire_switch_out_stage4[20]), .inData_21(wire_switch_out_stage4[21]), .inData_22(wire_switch_out_stage4[22]), .inData_23(wire_switch_out_stage4[23]), .inData_24(wire_switch_out_stage4[24]), .inData_25(wire_switch_out_stage4[25]), .inData_26(wire_switch_out_stage4[26]), .inData_27(wire_switch_out_stage4[27]), .inData_28(wire_switch_out_stage4[28]), .inData_29(wire_switch_out_stage4[29]), .inData_30(wire_switch_out_stage4[30]), .inData_31(wire_switch_out_stage4[31]), .inData_32(wire_switch_out_stage4[32]), .inData_33(wire_switch_out_stage4[33]), .inData_34(wire_switch_out_stage4[34]), .inData_35(wire_switch_out_stage4[35]), .inData_36(wire_switch_out_stage4[36]), .inData_37(wire_switch_out_stage4[37]), .inData_38(wire_switch_out_stage4[38]), .inData_39(wire_switch_out_stage4[39]), .inData_40(wire_switch_out_stage4[40]), .inData_41(wire_switch_out_stage4[41]), .inData_42(wire_switch_out_stage4[42]), .inData_43(wire_switch_out_stage4[43]), .inData_44(wire_switch_out_stage4[44]), .inData_45(wire_switch_out_stage4[45]), .inData_46(wire_switch_out_stage4[46]), .inData_47(wire_switch_out_stage4[47]), .inData_48(wire_switch_out_stage4[48]), .inData_49(wire_switch_out_stage4[49]), .inData_50(wire_switch_out_stage4[50]), .inData_51(wire_switch_out_stage4[51]), .inData_52(wire_switch_out_stage4[52]), .inData_53(wire_switch_out_stage4[53]), .inData_54(wire_switch_out_stage4[54]), .inData_55(wire_switch_out_stage4[55]), .inData_56(wire_switch_out_stage4[56]), .inData_57(wire_switch_out_stage4[57]), .inData_58(wire_switch_out_stage4[58]), .inData_59(wire_switch_out_stage4[59]), .inData_60(wire_switch_out_stage4[60]), .inData_61(wire_switch_out_stage4[61]), .inData_62(wire_switch_out_stage4[62]), .inData_63(wire_switch_out_stage4[63]), .inData_64(wire_switch_out_stage4[64]), .inData_65(wire_switch_out_stage4[65]), .inData_66(wire_switch_out_stage4[66]), .inData_67(wire_switch_out_stage4[67]), .inData_68(wire_switch_out_stage4[68]), .inData_69(wire_switch_out_stage4[69]), .inData_70(wire_switch_out_stage4[70]), .inData_71(wire_switch_out_stage4[71]), .inData_72(wire_switch_out_stage4[72]), .inData_73(wire_switch_out_stage4[73]), .inData_74(wire_switch_out_stage4[74]), .inData_75(wire_switch_out_stage4[75]), .inData_76(wire_switch_out_stage4[76]), .inData_77(wire_switch_out_stage4[77]), .inData_78(wire_switch_out_stage4[78]), .inData_79(wire_switch_out_stage4[79]), .inData_80(wire_switch_out_stage4[80]), .inData_81(wire_switch_out_stage4[81]), .inData_82(wire_switch_out_stage4[82]), .inData_83(wire_switch_out_stage4[83]), .inData_84(wire_switch_out_stage4[84]), .inData_85(wire_switch_out_stage4[85]), .inData_86(wire_switch_out_stage4[86]), .inData_87(wire_switch_out_stage4[87]), .inData_88(wire_switch_out_stage4[88]), .inData_89(wire_switch_out_stage4[89]), .inData_90(wire_switch_out_stage4[90]), .inData_91(wire_switch_out_stage4[91]), .inData_92(wire_switch_out_stage4[92]), .inData_93(wire_switch_out_stage4[93]), .inData_94(wire_switch_out_stage4[94]), .inData_95(wire_switch_out_stage4[95]), .inData_96(wire_switch_out_stage4[96]), .inData_97(wire_switch_out_stage4[97]), .inData_98(wire_switch_out_stage4[98]), .inData_99(wire_switch_out_stage4[99]), .inData_100(wire_switch_out_stage4[100]), .inData_101(wire_switch_out_stage4[101]), .inData_102(wire_switch_out_stage4[102]), .inData_103(wire_switch_out_stage4[103]), .inData_104(wire_switch_out_stage4[104]), .inData_105(wire_switch_out_stage4[105]), .inData_106(wire_switch_out_stage4[106]), .inData_107(wire_switch_out_stage4[107]), .inData_108(wire_switch_out_stage4[108]), .inData_109(wire_switch_out_stage4[109]), .inData_110(wire_switch_out_stage4[110]), .inData_111(wire_switch_out_stage4[111]), .inData_112(wire_switch_out_stage4[112]), .inData_113(wire_switch_out_stage4[113]), .inData_114(wire_switch_out_stage4[114]), .inData_115(wire_switch_out_stage4[115]), .inData_116(wire_switch_out_stage4[116]), .inData_117(wire_switch_out_stage4[117]), .inData_118(wire_switch_out_stage4[118]), .inData_119(wire_switch_out_stage4[119]), .inData_120(wire_switch_out_stage4[120]), .inData_121(wire_switch_out_stage4[121]), .inData_122(wire_switch_out_stage4[122]), .inData_123(wire_switch_out_stage4[123]), .inData_124(wire_switch_out_stage4[124]), .inData_125(wire_switch_out_stage4[125]), .inData_126(wire_switch_out_stage4[126]), .inData_127(wire_switch_out_stage4[127]), .inData_128(wire_switch_out_stage4[128]), .inData_129(wire_switch_out_stage4[129]), .inData_130(wire_switch_out_stage4[130]), .inData_131(wire_switch_out_stage4[131]), .inData_132(wire_switch_out_stage4[132]), .inData_133(wire_switch_out_stage4[133]), .inData_134(wire_switch_out_stage4[134]), .inData_135(wire_switch_out_stage4[135]), .inData_136(wire_switch_out_stage4[136]), .inData_137(wire_switch_out_stage4[137]), .inData_138(wire_switch_out_stage4[138]), .inData_139(wire_switch_out_stage4[139]), .inData_140(wire_switch_out_stage4[140]), .inData_141(wire_switch_out_stage4[141]), .inData_142(wire_switch_out_stage4[142]), .inData_143(wire_switch_out_stage4[143]), .inData_144(wire_switch_out_stage4[144]), .inData_145(wire_switch_out_stage4[145]), .inData_146(wire_switch_out_stage4[146]), .inData_147(wire_switch_out_stage4[147]), .inData_148(wire_switch_out_stage4[148]), .inData_149(wire_switch_out_stage4[149]), .inData_150(wire_switch_out_stage4[150]), .inData_151(wire_switch_out_stage4[151]), .inData_152(wire_switch_out_stage4[152]), .inData_153(wire_switch_out_stage4[153]), .inData_154(wire_switch_out_stage4[154]), .inData_155(wire_switch_out_stage4[155]), .inData_156(wire_switch_out_stage4[156]), .inData_157(wire_switch_out_stage4[157]), .inData_158(wire_switch_out_stage4[158]), .inData_159(wire_switch_out_stage4[159]), .inData_160(wire_switch_out_stage4[160]), .inData_161(wire_switch_out_stage4[161]), .inData_162(wire_switch_out_stage4[162]), .inData_163(wire_switch_out_stage4[163]), .inData_164(wire_switch_out_stage4[164]), .inData_165(wire_switch_out_stage4[165]), .inData_166(wire_switch_out_stage4[166]), .inData_167(wire_switch_out_stage4[167]), .inData_168(wire_switch_out_stage4[168]), .inData_169(wire_switch_out_stage4[169]), .inData_170(wire_switch_out_stage4[170]), .inData_171(wire_switch_out_stage4[171]), .inData_172(wire_switch_out_stage4[172]), .inData_173(wire_switch_out_stage4[173]), .inData_174(wire_switch_out_stage4[174]), .inData_175(wire_switch_out_stage4[175]), .inData_176(wire_switch_out_stage4[176]), .inData_177(wire_switch_out_stage4[177]), .inData_178(wire_switch_out_stage4[178]), .inData_179(wire_switch_out_stage4[179]), .inData_180(wire_switch_out_stage4[180]), .inData_181(wire_switch_out_stage4[181]), .inData_182(wire_switch_out_stage4[182]), .inData_183(wire_switch_out_stage4[183]), .inData_184(wire_switch_out_stage4[184]), .inData_185(wire_switch_out_stage4[185]), .inData_186(wire_switch_out_stage4[186]), .inData_187(wire_switch_out_stage4[187]), .inData_188(wire_switch_out_stage4[188]), .inData_189(wire_switch_out_stage4[189]), .inData_190(wire_switch_out_stage4[190]), .inData_191(wire_switch_out_stage4[191]), .inData_192(wire_switch_out_stage4[192]), .inData_193(wire_switch_out_stage4[193]), .inData_194(wire_switch_out_stage4[194]), .inData_195(wire_switch_out_stage4[195]), .inData_196(wire_switch_out_stage4[196]), .inData_197(wire_switch_out_stage4[197]), .inData_198(wire_switch_out_stage4[198]), .inData_199(wire_switch_out_stage4[199]), .inData_200(wire_switch_out_stage4[200]), .inData_201(wire_switch_out_stage4[201]), .inData_202(wire_switch_out_stage4[202]), .inData_203(wire_switch_out_stage4[203]), .inData_204(wire_switch_out_stage4[204]), .inData_205(wire_switch_out_stage4[205]), .inData_206(wire_switch_out_stage4[206]), .inData_207(wire_switch_out_stage4[207]), .inData_208(wire_switch_out_stage4[208]), .inData_209(wire_switch_out_stage4[209]), .inData_210(wire_switch_out_stage4[210]), .inData_211(wire_switch_out_stage4[211]), .inData_212(wire_switch_out_stage4[212]), .inData_213(wire_switch_out_stage4[213]), .inData_214(wire_switch_out_stage4[214]), .inData_215(wire_switch_out_stage4[215]), .inData_216(wire_switch_out_stage4[216]), .inData_217(wire_switch_out_stage4[217]), .inData_218(wire_switch_out_stage4[218]), .inData_219(wire_switch_out_stage4[219]), .inData_220(wire_switch_out_stage4[220]), .inData_221(wire_switch_out_stage4[221]), .inData_222(wire_switch_out_stage4[222]), .inData_223(wire_switch_out_stage4[223]), .inData_224(wire_switch_out_stage4[224]), .inData_225(wire_switch_out_stage4[225]), .inData_226(wire_switch_out_stage4[226]), .inData_227(wire_switch_out_stage4[227]), .inData_228(wire_switch_out_stage4[228]), .inData_229(wire_switch_out_stage4[229]), .inData_230(wire_switch_out_stage4[230]), .inData_231(wire_switch_out_stage4[231]), .inData_232(wire_switch_out_stage4[232]), .inData_233(wire_switch_out_stage4[233]), .inData_234(wire_switch_out_stage4[234]), .inData_235(wire_switch_out_stage4[235]), .inData_236(wire_switch_out_stage4[236]), .inData_237(wire_switch_out_stage4[237]), .inData_238(wire_switch_out_stage4[238]), .inData_239(wire_switch_out_stage4[239]), .inData_240(wire_switch_out_stage4[240]), .inData_241(wire_switch_out_stage4[241]), .inData_242(wire_switch_out_stage4[242]), .inData_243(wire_switch_out_stage4[243]), .inData_244(wire_switch_out_stage4[244]), .inData_245(wire_switch_out_stage4[245]), .inData_246(wire_switch_out_stage4[246]), .inData_247(wire_switch_out_stage4[247]), .inData_248(wire_switch_out_stage4[248]), .inData_249(wire_switch_out_stage4[249]), .inData_250(wire_switch_out_stage4[250]), .inData_251(wire_switch_out_stage4[251]), .inData_252(wire_switch_out_stage4[252]), .inData_253(wire_switch_out_stage4[253]), .inData_254(wire_switch_out_stage4[254]), .inData_255(wire_switch_out_stage4[255]), 
        .outData_0(wire_switch_in_stage3[0]), .outData_1(wire_switch_in_stage3[1]), .outData_2(wire_switch_in_stage3[2]), .outData_3(wire_switch_in_stage3[3]), .outData_4(wire_switch_in_stage3[4]), .outData_5(wire_switch_in_stage3[5]), .outData_6(wire_switch_in_stage3[6]), .outData_7(wire_switch_in_stage3[7]), .outData_8(wire_switch_in_stage3[8]), .outData_9(wire_switch_in_stage3[9]), .outData_10(wire_switch_in_stage3[10]), .outData_11(wire_switch_in_stage3[11]), .outData_12(wire_switch_in_stage3[12]), .outData_13(wire_switch_in_stage3[13]), .outData_14(wire_switch_in_stage3[14]), .outData_15(wire_switch_in_stage3[15]), .outData_16(wire_switch_in_stage3[16]), .outData_17(wire_switch_in_stage3[17]), .outData_18(wire_switch_in_stage3[18]), .outData_19(wire_switch_in_stage3[19]), .outData_20(wire_switch_in_stage3[20]), .outData_21(wire_switch_in_stage3[21]), .outData_22(wire_switch_in_stage3[22]), .outData_23(wire_switch_in_stage3[23]), .outData_24(wire_switch_in_stage3[24]), .outData_25(wire_switch_in_stage3[25]), .outData_26(wire_switch_in_stage3[26]), .outData_27(wire_switch_in_stage3[27]), .outData_28(wire_switch_in_stage3[28]), .outData_29(wire_switch_in_stage3[29]), .outData_30(wire_switch_in_stage3[30]), .outData_31(wire_switch_in_stage3[31]), .outData_32(wire_switch_in_stage3[32]), .outData_33(wire_switch_in_stage3[33]), .outData_34(wire_switch_in_stage3[34]), .outData_35(wire_switch_in_stage3[35]), .outData_36(wire_switch_in_stage3[36]), .outData_37(wire_switch_in_stage3[37]), .outData_38(wire_switch_in_stage3[38]), .outData_39(wire_switch_in_stage3[39]), .outData_40(wire_switch_in_stage3[40]), .outData_41(wire_switch_in_stage3[41]), .outData_42(wire_switch_in_stage3[42]), .outData_43(wire_switch_in_stage3[43]), .outData_44(wire_switch_in_stage3[44]), .outData_45(wire_switch_in_stage3[45]), .outData_46(wire_switch_in_stage3[46]), .outData_47(wire_switch_in_stage3[47]), .outData_48(wire_switch_in_stage3[48]), .outData_49(wire_switch_in_stage3[49]), .outData_50(wire_switch_in_stage3[50]), .outData_51(wire_switch_in_stage3[51]), .outData_52(wire_switch_in_stage3[52]), .outData_53(wire_switch_in_stage3[53]), .outData_54(wire_switch_in_stage3[54]), .outData_55(wire_switch_in_stage3[55]), .outData_56(wire_switch_in_stage3[56]), .outData_57(wire_switch_in_stage3[57]), .outData_58(wire_switch_in_stage3[58]), .outData_59(wire_switch_in_stage3[59]), .outData_60(wire_switch_in_stage3[60]), .outData_61(wire_switch_in_stage3[61]), .outData_62(wire_switch_in_stage3[62]), .outData_63(wire_switch_in_stage3[63]), .outData_64(wire_switch_in_stage3[64]), .outData_65(wire_switch_in_stage3[65]), .outData_66(wire_switch_in_stage3[66]), .outData_67(wire_switch_in_stage3[67]), .outData_68(wire_switch_in_stage3[68]), .outData_69(wire_switch_in_stage3[69]), .outData_70(wire_switch_in_stage3[70]), .outData_71(wire_switch_in_stage3[71]), .outData_72(wire_switch_in_stage3[72]), .outData_73(wire_switch_in_stage3[73]), .outData_74(wire_switch_in_stage3[74]), .outData_75(wire_switch_in_stage3[75]), .outData_76(wire_switch_in_stage3[76]), .outData_77(wire_switch_in_stage3[77]), .outData_78(wire_switch_in_stage3[78]), .outData_79(wire_switch_in_stage3[79]), .outData_80(wire_switch_in_stage3[80]), .outData_81(wire_switch_in_stage3[81]), .outData_82(wire_switch_in_stage3[82]), .outData_83(wire_switch_in_stage3[83]), .outData_84(wire_switch_in_stage3[84]), .outData_85(wire_switch_in_stage3[85]), .outData_86(wire_switch_in_stage3[86]), .outData_87(wire_switch_in_stage3[87]), .outData_88(wire_switch_in_stage3[88]), .outData_89(wire_switch_in_stage3[89]), .outData_90(wire_switch_in_stage3[90]), .outData_91(wire_switch_in_stage3[91]), .outData_92(wire_switch_in_stage3[92]), .outData_93(wire_switch_in_stage3[93]), .outData_94(wire_switch_in_stage3[94]), .outData_95(wire_switch_in_stage3[95]), .outData_96(wire_switch_in_stage3[96]), .outData_97(wire_switch_in_stage3[97]), .outData_98(wire_switch_in_stage3[98]), .outData_99(wire_switch_in_stage3[99]), .outData_100(wire_switch_in_stage3[100]), .outData_101(wire_switch_in_stage3[101]), .outData_102(wire_switch_in_stage3[102]), .outData_103(wire_switch_in_stage3[103]), .outData_104(wire_switch_in_stage3[104]), .outData_105(wire_switch_in_stage3[105]), .outData_106(wire_switch_in_stage3[106]), .outData_107(wire_switch_in_stage3[107]), .outData_108(wire_switch_in_stage3[108]), .outData_109(wire_switch_in_stage3[109]), .outData_110(wire_switch_in_stage3[110]), .outData_111(wire_switch_in_stage3[111]), .outData_112(wire_switch_in_stage3[112]), .outData_113(wire_switch_in_stage3[113]), .outData_114(wire_switch_in_stage3[114]), .outData_115(wire_switch_in_stage3[115]), .outData_116(wire_switch_in_stage3[116]), .outData_117(wire_switch_in_stage3[117]), .outData_118(wire_switch_in_stage3[118]), .outData_119(wire_switch_in_stage3[119]), .outData_120(wire_switch_in_stage3[120]), .outData_121(wire_switch_in_stage3[121]), .outData_122(wire_switch_in_stage3[122]), .outData_123(wire_switch_in_stage3[123]), .outData_124(wire_switch_in_stage3[124]), .outData_125(wire_switch_in_stage3[125]), .outData_126(wire_switch_in_stage3[126]), .outData_127(wire_switch_in_stage3[127]), .outData_128(wire_switch_in_stage3[128]), .outData_129(wire_switch_in_stage3[129]), .outData_130(wire_switch_in_stage3[130]), .outData_131(wire_switch_in_stage3[131]), .outData_132(wire_switch_in_stage3[132]), .outData_133(wire_switch_in_stage3[133]), .outData_134(wire_switch_in_stage3[134]), .outData_135(wire_switch_in_stage3[135]), .outData_136(wire_switch_in_stage3[136]), .outData_137(wire_switch_in_stage3[137]), .outData_138(wire_switch_in_stage3[138]), .outData_139(wire_switch_in_stage3[139]), .outData_140(wire_switch_in_stage3[140]), .outData_141(wire_switch_in_stage3[141]), .outData_142(wire_switch_in_stage3[142]), .outData_143(wire_switch_in_stage3[143]), .outData_144(wire_switch_in_stage3[144]), .outData_145(wire_switch_in_stage3[145]), .outData_146(wire_switch_in_stage3[146]), .outData_147(wire_switch_in_stage3[147]), .outData_148(wire_switch_in_stage3[148]), .outData_149(wire_switch_in_stage3[149]), .outData_150(wire_switch_in_stage3[150]), .outData_151(wire_switch_in_stage3[151]), .outData_152(wire_switch_in_stage3[152]), .outData_153(wire_switch_in_stage3[153]), .outData_154(wire_switch_in_stage3[154]), .outData_155(wire_switch_in_stage3[155]), .outData_156(wire_switch_in_stage3[156]), .outData_157(wire_switch_in_stage3[157]), .outData_158(wire_switch_in_stage3[158]), .outData_159(wire_switch_in_stage3[159]), .outData_160(wire_switch_in_stage3[160]), .outData_161(wire_switch_in_stage3[161]), .outData_162(wire_switch_in_stage3[162]), .outData_163(wire_switch_in_stage3[163]), .outData_164(wire_switch_in_stage3[164]), .outData_165(wire_switch_in_stage3[165]), .outData_166(wire_switch_in_stage3[166]), .outData_167(wire_switch_in_stage3[167]), .outData_168(wire_switch_in_stage3[168]), .outData_169(wire_switch_in_stage3[169]), .outData_170(wire_switch_in_stage3[170]), .outData_171(wire_switch_in_stage3[171]), .outData_172(wire_switch_in_stage3[172]), .outData_173(wire_switch_in_stage3[173]), .outData_174(wire_switch_in_stage3[174]), .outData_175(wire_switch_in_stage3[175]), .outData_176(wire_switch_in_stage3[176]), .outData_177(wire_switch_in_stage3[177]), .outData_178(wire_switch_in_stage3[178]), .outData_179(wire_switch_in_stage3[179]), .outData_180(wire_switch_in_stage3[180]), .outData_181(wire_switch_in_stage3[181]), .outData_182(wire_switch_in_stage3[182]), .outData_183(wire_switch_in_stage3[183]), .outData_184(wire_switch_in_stage3[184]), .outData_185(wire_switch_in_stage3[185]), .outData_186(wire_switch_in_stage3[186]), .outData_187(wire_switch_in_stage3[187]), .outData_188(wire_switch_in_stage3[188]), .outData_189(wire_switch_in_stage3[189]), .outData_190(wire_switch_in_stage3[190]), .outData_191(wire_switch_in_stage3[191]), .outData_192(wire_switch_in_stage3[192]), .outData_193(wire_switch_in_stage3[193]), .outData_194(wire_switch_in_stage3[194]), .outData_195(wire_switch_in_stage3[195]), .outData_196(wire_switch_in_stage3[196]), .outData_197(wire_switch_in_stage3[197]), .outData_198(wire_switch_in_stage3[198]), .outData_199(wire_switch_in_stage3[199]), .outData_200(wire_switch_in_stage3[200]), .outData_201(wire_switch_in_stage3[201]), .outData_202(wire_switch_in_stage3[202]), .outData_203(wire_switch_in_stage3[203]), .outData_204(wire_switch_in_stage3[204]), .outData_205(wire_switch_in_stage3[205]), .outData_206(wire_switch_in_stage3[206]), .outData_207(wire_switch_in_stage3[207]), .outData_208(wire_switch_in_stage3[208]), .outData_209(wire_switch_in_stage3[209]), .outData_210(wire_switch_in_stage3[210]), .outData_211(wire_switch_in_stage3[211]), .outData_212(wire_switch_in_stage3[212]), .outData_213(wire_switch_in_stage3[213]), .outData_214(wire_switch_in_stage3[214]), .outData_215(wire_switch_in_stage3[215]), .outData_216(wire_switch_in_stage3[216]), .outData_217(wire_switch_in_stage3[217]), .outData_218(wire_switch_in_stage3[218]), .outData_219(wire_switch_in_stage3[219]), .outData_220(wire_switch_in_stage3[220]), .outData_221(wire_switch_in_stage3[221]), .outData_222(wire_switch_in_stage3[222]), .outData_223(wire_switch_in_stage3[223]), .outData_224(wire_switch_in_stage3[224]), .outData_225(wire_switch_in_stage3[225]), .outData_226(wire_switch_in_stage3[226]), .outData_227(wire_switch_in_stage3[227]), .outData_228(wire_switch_in_stage3[228]), .outData_229(wire_switch_in_stage3[229]), .outData_230(wire_switch_in_stage3[230]), .outData_231(wire_switch_in_stage3[231]), .outData_232(wire_switch_in_stage3[232]), .outData_233(wire_switch_in_stage3[233]), .outData_234(wire_switch_in_stage3[234]), .outData_235(wire_switch_in_stage3[235]), .outData_236(wire_switch_in_stage3[236]), .outData_237(wire_switch_in_stage3[237]), .outData_238(wire_switch_in_stage3[238]), .outData_239(wire_switch_in_stage3[239]), .outData_240(wire_switch_in_stage3[240]), .outData_241(wire_switch_in_stage3[241]), .outData_242(wire_switch_in_stage3[242]), .outData_243(wire_switch_in_stage3[243]), .outData_244(wire_switch_in_stage3[244]), .outData_245(wire_switch_in_stage3[245]), .outData_246(wire_switch_in_stage3[246]), .outData_247(wire_switch_in_stage3[247]), .outData_248(wire_switch_in_stage3[248]), .outData_249(wire_switch_in_stage3[249]), .outData_250(wire_switch_in_stage3[250]), .outData_251(wire_switch_in_stage3[251]), .outData_252(wire_switch_in_stage3[252]), .outData_253(wire_switch_in_stage3[253]), .outData_254(wire_switch_in_stage3[254]), .outData_255(wire_switch_in_stage3[255]), 
        .in_start(in_start_stage3), .out_start(con_in_start_stage3), .clk(clk), .rst(rst)); 

  
  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[0] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[1] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[2] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[3] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[4] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[5] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[6] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[7] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[8] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[9] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[10] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[11] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[12] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[13] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[14] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[15] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[16] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[17] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[18] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[19] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[20] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[21] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[22] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[23] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[24] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[25] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[26] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[27] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[28] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[29] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[30] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[31] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[32] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[33] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[34] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[35] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[36] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[37] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[38] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[39] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[40] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[41] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[42] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[43] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[44] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[45] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[46] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[47] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[48] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[49] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[50] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[51] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[52] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[53] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[54] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[55] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[56] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[57] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[58] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[59] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[60] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[61] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[62] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[63] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[64] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[65] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[66] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[67] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[68] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[69] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[70] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[71] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[72] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[73] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[74] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[75] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[76] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[77] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[78] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[79] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[80] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[81] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[82] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[83] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[84] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[85] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[86] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[87] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[88] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[89] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[90] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[91] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[92] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[93] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[94] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[95] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[96] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[97] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[98] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[99] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[100] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[101] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[102] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[103] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[104] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[105] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[106] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[107] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[108] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[109] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[110] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[111] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[112] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[113] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[114] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[115] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[116] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[117] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[118] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[119] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[120] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[121] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[122] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[123] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[124] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[125] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[126] <= counter_w[4]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage3[127] <= counter_w[4]; 
  end                            

  wire [DATA_WIDTH-1:0] wire_switch_in_stage2[255:0];
  wire [DATA_WIDTH-1:0] wire_switch_out_stage2[255:0];
  reg [127:0] wire_ctrl_stage2;

  switches_stage_st2_0_R switch_stage_2(
        .inData_0(wire_switch_in_stage2[0]), .inData_1(wire_switch_in_stage2[1]), .inData_2(wire_switch_in_stage2[2]), .inData_3(wire_switch_in_stage2[3]), .inData_4(wire_switch_in_stage2[4]), .inData_5(wire_switch_in_stage2[5]), .inData_6(wire_switch_in_stage2[6]), .inData_7(wire_switch_in_stage2[7]), .inData_8(wire_switch_in_stage2[8]), .inData_9(wire_switch_in_stage2[9]), .inData_10(wire_switch_in_stage2[10]), .inData_11(wire_switch_in_stage2[11]), .inData_12(wire_switch_in_stage2[12]), .inData_13(wire_switch_in_stage2[13]), .inData_14(wire_switch_in_stage2[14]), .inData_15(wire_switch_in_stage2[15]), .inData_16(wire_switch_in_stage2[16]), .inData_17(wire_switch_in_stage2[17]), .inData_18(wire_switch_in_stage2[18]), .inData_19(wire_switch_in_stage2[19]), .inData_20(wire_switch_in_stage2[20]), .inData_21(wire_switch_in_stage2[21]), .inData_22(wire_switch_in_stage2[22]), .inData_23(wire_switch_in_stage2[23]), .inData_24(wire_switch_in_stage2[24]), .inData_25(wire_switch_in_stage2[25]), .inData_26(wire_switch_in_stage2[26]), .inData_27(wire_switch_in_stage2[27]), .inData_28(wire_switch_in_stage2[28]), .inData_29(wire_switch_in_stage2[29]), .inData_30(wire_switch_in_stage2[30]), .inData_31(wire_switch_in_stage2[31]), .inData_32(wire_switch_in_stage2[32]), .inData_33(wire_switch_in_stage2[33]), .inData_34(wire_switch_in_stage2[34]), .inData_35(wire_switch_in_stage2[35]), .inData_36(wire_switch_in_stage2[36]), .inData_37(wire_switch_in_stage2[37]), .inData_38(wire_switch_in_stage2[38]), .inData_39(wire_switch_in_stage2[39]), .inData_40(wire_switch_in_stage2[40]), .inData_41(wire_switch_in_stage2[41]), .inData_42(wire_switch_in_stage2[42]), .inData_43(wire_switch_in_stage2[43]), .inData_44(wire_switch_in_stage2[44]), .inData_45(wire_switch_in_stage2[45]), .inData_46(wire_switch_in_stage2[46]), .inData_47(wire_switch_in_stage2[47]), .inData_48(wire_switch_in_stage2[48]), .inData_49(wire_switch_in_stage2[49]), .inData_50(wire_switch_in_stage2[50]), .inData_51(wire_switch_in_stage2[51]), .inData_52(wire_switch_in_stage2[52]), .inData_53(wire_switch_in_stage2[53]), .inData_54(wire_switch_in_stage2[54]), .inData_55(wire_switch_in_stage2[55]), .inData_56(wire_switch_in_stage2[56]), .inData_57(wire_switch_in_stage2[57]), .inData_58(wire_switch_in_stage2[58]), .inData_59(wire_switch_in_stage2[59]), .inData_60(wire_switch_in_stage2[60]), .inData_61(wire_switch_in_stage2[61]), .inData_62(wire_switch_in_stage2[62]), .inData_63(wire_switch_in_stage2[63]), .inData_64(wire_switch_in_stage2[64]), .inData_65(wire_switch_in_stage2[65]), .inData_66(wire_switch_in_stage2[66]), .inData_67(wire_switch_in_stage2[67]), .inData_68(wire_switch_in_stage2[68]), .inData_69(wire_switch_in_stage2[69]), .inData_70(wire_switch_in_stage2[70]), .inData_71(wire_switch_in_stage2[71]), .inData_72(wire_switch_in_stage2[72]), .inData_73(wire_switch_in_stage2[73]), .inData_74(wire_switch_in_stage2[74]), .inData_75(wire_switch_in_stage2[75]), .inData_76(wire_switch_in_stage2[76]), .inData_77(wire_switch_in_stage2[77]), .inData_78(wire_switch_in_stage2[78]), .inData_79(wire_switch_in_stage2[79]), .inData_80(wire_switch_in_stage2[80]), .inData_81(wire_switch_in_stage2[81]), .inData_82(wire_switch_in_stage2[82]), .inData_83(wire_switch_in_stage2[83]), .inData_84(wire_switch_in_stage2[84]), .inData_85(wire_switch_in_stage2[85]), .inData_86(wire_switch_in_stage2[86]), .inData_87(wire_switch_in_stage2[87]), .inData_88(wire_switch_in_stage2[88]), .inData_89(wire_switch_in_stage2[89]), .inData_90(wire_switch_in_stage2[90]), .inData_91(wire_switch_in_stage2[91]), .inData_92(wire_switch_in_stage2[92]), .inData_93(wire_switch_in_stage2[93]), .inData_94(wire_switch_in_stage2[94]), .inData_95(wire_switch_in_stage2[95]), .inData_96(wire_switch_in_stage2[96]), .inData_97(wire_switch_in_stage2[97]), .inData_98(wire_switch_in_stage2[98]), .inData_99(wire_switch_in_stage2[99]), .inData_100(wire_switch_in_stage2[100]), .inData_101(wire_switch_in_stage2[101]), .inData_102(wire_switch_in_stage2[102]), .inData_103(wire_switch_in_stage2[103]), .inData_104(wire_switch_in_stage2[104]), .inData_105(wire_switch_in_stage2[105]), .inData_106(wire_switch_in_stage2[106]), .inData_107(wire_switch_in_stage2[107]), .inData_108(wire_switch_in_stage2[108]), .inData_109(wire_switch_in_stage2[109]), .inData_110(wire_switch_in_stage2[110]), .inData_111(wire_switch_in_stage2[111]), .inData_112(wire_switch_in_stage2[112]), .inData_113(wire_switch_in_stage2[113]), .inData_114(wire_switch_in_stage2[114]), .inData_115(wire_switch_in_stage2[115]), .inData_116(wire_switch_in_stage2[116]), .inData_117(wire_switch_in_stage2[117]), .inData_118(wire_switch_in_stage2[118]), .inData_119(wire_switch_in_stage2[119]), .inData_120(wire_switch_in_stage2[120]), .inData_121(wire_switch_in_stage2[121]), .inData_122(wire_switch_in_stage2[122]), .inData_123(wire_switch_in_stage2[123]), .inData_124(wire_switch_in_stage2[124]), .inData_125(wire_switch_in_stage2[125]), .inData_126(wire_switch_in_stage2[126]), .inData_127(wire_switch_in_stage2[127]), .inData_128(wire_switch_in_stage2[128]), .inData_129(wire_switch_in_stage2[129]), .inData_130(wire_switch_in_stage2[130]), .inData_131(wire_switch_in_stage2[131]), .inData_132(wire_switch_in_stage2[132]), .inData_133(wire_switch_in_stage2[133]), .inData_134(wire_switch_in_stage2[134]), .inData_135(wire_switch_in_stage2[135]), .inData_136(wire_switch_in_stage2[136]), .inData_137(wire_switch_in_stage2[137]), .inData_138(wire_switch_in_stage2[138]), .inData_139(wire_switch_in_stage2[139]), .inData_140(wire_switch_in_stage2[140]), .inData_141(wire_switch_in_stage2[141]), .inData_142(wire_switch_in_stage2[142]), .inData_143(wire_switch_in_stage2[143]), .inData_144(wire_switch_in_stage2[144]), .inData_145(wire_switch_in_stage2[145]), .inData_146(wire_switch_in_stage2[146]), .inData_147(wire_switch_in_stage2[147]), .inData_148(wire_switch_in_stage2[148]), .inData_149(wire_switch_in_stage2[149]), .inData_150(wire_switch_in_stage2[150]), .inData_151(wire_switch_in_stage2[151]), .inData_152(wire_switch_in_stage2[152]), .inData_153(wire_switch_in_stage2[153]), .inData_154(wire_switch_in_stage2[154]), .inData_155(wire_switch_in_stage2[155]), .inData_156(wire_switch_in_stage2[156]), .inData_157(wire_switch_in_stage2[157]), .inData_158(wire_switch_in_stage2[158]), .inData_159(wire_switch_in_stage2[159]), .inData_160(wire_switch_in_stage2[160]), .inData_161(wire_switch_in_stage2[161]), .inData_162(wire_switch_in_stage2[162]), .inData_163(wire_switch_in_stage2[163]), .inData_164(wire_switch_in_stage2[164]), .inData_165(wire_switch_in_stage2[165]), .inData_166(wire_switch_in_stage2[166]), .inData_167(wire_switch_in_stage2[167]), .inData_168(wire_switch_in_stage2[168]), .inData_169(wire_switch_in_stage2[169]), .inData_170(wire_switch_in_stage2[170]), .inData_171(wire_switch_in_stage2[171]), .inData_172(wire_switch_in_stage2[172]), .inData_173(wire_switch_in_stage2[173]), .inData_174(wire_switch_in_stage2[174]), .inData_175(wire_switch_in_stage2[175]), .inData_176(wire_switch_in_stage2[176]), .inData_177(wire_switch_in_stage2[177]), .inData_178(wire_switch_in_stage2[178]), .inData_179(wire_switch_in_stage2[179]), .inData_180(wire_switch_in_stage2[180]), .inData_181(wire_switch_in_stage2[181]), .inData_182(wire_switch_in_stage2[182]), .inData_183(wire_switch_in_stage2[183]), .inData_184(wire_switch_in_stage2[184]), .inData_185(wire_switch_in_stage2[185]), .inData_186(wire_switch_in_stage2[186]), .inData_187(wire_switch_in_stage2[187]), .inData_188(wire_switch_in_stage2[188]), .inData_189(wire_switch_in_stage2[189]), .inData_190(wire_switch_in_stage2[190]), .inData_191(wire_switch_in_stage2[191]), .inData_192(wire_switch_in_stage2[192]), .inData_193(wire_switch_in_stage2[193]), .inData_194(wire_switch_in_stage2[194]), .inData_195(wire_switch_in_stage2[195]), .inData_196(wire_switch_in_stage2[196]), .inData_197(wire_switch_in_stage2[197]), .inData_198(wire_switch_in_stage2[198]), .inData_199(wire_switch_in_stage2[199]), .inData_200(wire_switch_in_stage2[200]), .inData_201(wire_switch_in_stage2[201]), .inData_202(wire_switch_in_stage2[202]), .inData_203(wire_switch_in_stage2[203]), .inData_204(wire_switch_in_stage2[204]), .inData_205(wire_switch_in_stage2[205]), .inData_206(wire_switch_in_stage2[206]), .inData_207(wire_switch_in_stage2[207]), .inData_208(wire_switch_in_stage2[208]), .inData_209(wire_switch_in_stage2[209]), .inData_210(wire_switch_in_stage2[210]), .inData_211(wire_switch_in_stage2[211]), .inData_212(wire_switch_in_stage2[212]), .inData_213(wire_switch_in_stage2[213]), .inData_214(wire_switch_in_stage2[214]), .inData_215(wire_switch_in_stage2[215]), .inData_216(wire_switch_in_stage2[216]), .inData_217(wire_switch_in_stage2[217]), .inData_218(wire_switch_in_stage2[218]), .inData_219(wire_switch_in_stage2[219]), .inData_220(wire_switch_in_stage2[220]), .inData_221(wire_switch_in_stage2[221]), .inData_222(wire_switch_in_stage2[222]), .inData_223(wire_switch_in_stage2[223]), .inData_224(wire_switch_in_stage2[224]), .inData_225(wire_switch_in_stage2[225]), .inData_226(wire_switch_in_stage2[226]), .inData_227(wire_switch_in_stage2[227]), .inData_228(wire_switch_in_stage2[228]), .inData_229(wire_switch_in_stage2[229]), .inData_230(wire_switch_in_stage2[230]), .inData_231(wire_switch_in_stage2[231]), .inData_232(wire_switch_in_stage2[232]), .inData_233(wire_switch_in_stage2[233]), .inData_234(wire_switch_in_stage2[234]), .inData_235(wire_switch_in_stage2[235]), .inData_236(wire_switch_in_stage2[236]), .inData_237(wire_switch_in_stage2[237]), .inData_238(wire_switch_in_stage2[238]), .inData_239(wire_switch_in_stage2[239]), .inData_240(wire_switch_in_stage2[240]), .inData_241(wire_switch_in_stage2[241]), .inData_242(wire_switch_in_stage2[242]), .inData_243(wire_switch_in_stage2[243]), .inData_244(wire_switch_in_stage2[244]), .inData_245(wire_switch_in_stage2[245]), .inData_246(wire_switch_in_stage2[246]), .inData_247(wire_switch_in_stage2[247]), .inData_248(wire_switch_in_stage2[248]), .inData_249(wire_switch_in_stage2[249]), .inData_250(wire_switch_in_stage2[250]), .inData_251(wire_switch_in_stage2[251]), .inData_252(wire_switch_in_stage2[252]), .inData_253(wire_switch_in_stage2[253]), .inData_254(wire_switch_in_stage2[254]), .inData_255(wire_switch_in_stage2[255]), 
        .outData_0(wire_switch_out_stage2[0]), .outData_1(wire_switch_out_stage2[1]), .outData_2(wire_switch_out_stage2[2]), .outData_3(wire_switch_out_stage2[3]), .outData_4(wire_switch_out_stage2[4]), .outData_5(wire_switch_out_stage2[5]), .outData_6(wire_switch_out_stage2[6]), .outData_7(wire_switch_out_stage2[7]), .outData_8(wire_switch_out_stage2[8]), .outData_9(wire_switch_out_stage2[9]), .outData_10(wire_switch_out_stage2[10]), .outData_11(wire_switch_out_stage2[11]), .outData_12(wire_switch_out_stage2[12]), .outData_13(wire_switch_out_stage2[13]), .outData_14(wire_switch_out_stage2[14]), .outData_15(wire_switch_out_stage2[15]), .outData_16(wire_switch_out_stage2[16]), .outData_17(wire_switch_out_stage2[17]), .outData_18(wire_switch_out_stage2[18]), .outData_19(wire_switch_out_stage2[19]), .outData_20(wire_switch_out_stage2[20]), .outData_21(wire_switch_out_stage2[21]), .outData_22(wire_switch_out_stage2[22]), .outData_23(wire_switch_out_stage2[23]), .outData_24(wire_switch_out_stage2[24]), .outData_25(wire_switch_out_stage2[25]), .outData_26(wire_switch_out_stage2[26]), .outData_27(wire_switch_out_stage2[27]), .outData_28(wire_switch_out_stage2[28]), .outData_29(wire_switch_out_stage2[29]), .outData_30(wire_switch_out_stage2[30]), .outData_31(wire_switch_out_stage2[31]), .outData_32(wire_switch_out_stage2[32]), .outData_33(wire_switch_out_stage2[33]), .outData_34(wire_switch_out_stage2[34]), .outData_35(wire_switch_out_stage2[35]), .outData_36(wire_switch_out_stage2[36]), .outData_37(wire_switch_out_stage2[37]), .outData_38(wire_switch_out_stage2[38]), .outData_39(wire_switch_out_stage2[39]), .outData_40(wire_switch_out_stage2[40]), .outData_41(wire_switch_out_stage2[41]), .outData_42(wire_switch_out_stage2[42]), .outData_43(wire_switch_out_stage2[43]), .outData_44(wire_switch_out_stage2[44]), .outData_45(wire_switch_out_stage2[45]), .outData_46(wire_switch_out_stage2[46]), .outData_47(wire_switch_out_stage2[47]), .outData_48(wire_switch_out_stage2[48]), .outData_49(wire_switch_out_stage2[49]), .outData_50(wire_switch_out_stage2[50]), .outData_51(wire_switch_out_stage2[51]), .outData_52(wire_switch_out_stage2[52]), .outData_53(wire_switch_out_stage2[53]), .outData_54(wire_switch_out_stage2[54]), .outData_55(wire_switch_out_stage2[55]), .outData_56(wire_switch_out_stage2[56]), .outData_57(wire_switch_out_stage2[57]), .outData_58(wire_switch_out_stage2[58]), .outData_59(wire_switch_out_stage2[59]), .outData_60(wire_switch_out_stage2[60]), .outData_61(wire_switch_out_stage2[61]), .outData_62(wire_switch_out_stage2[62]), .outData_63(wire_switch_out_stage2[63]), .outData_64(wire_switch_out_stage2[64]), .outData_65(wire_switch_out_stage2[65]), .outData_66(wire_switch_out_stage2[66]), .outData_67(wire_switch_out_stage2[67]), .outData_68(wire_switch_out_stage2[68]), .outData_69(wire_switch_out_stage2[69]), .outData_70(wire_switch_out_stage2[70]), .outData_71(wire_switch_out_stage2[71]), .outData_72(wire_switch_out_stage2[72]), .outData_73(wire_switch_out_stage2[73]), .outData_74(wire_switch_out_stage2[74]), .outData_75(wire_switch_out_stage2[75]), .outData_76(wire_switch_out_stage2[76]), .outData_77(wire_switch_out_stage2[77]), .outData_78(wire_switch_out_stage2[78]), .outData_79(wire_switch_out_stage2[79]), .outData_80(wire_switch_out_stage2[80]), .outData_81(wire_switch_out_stage2[81]), .outData_82(wire_switch_out_stage2[82]), .outData_83(wire_switch_out_stage2[83]), .outData_84(wire_switch_out_stage2[84]), .outData_85(wire_switch_out_stage2[85]), .outData_86(wire_switch_out_stage2[86]), .outData_87(wire_switch_out_stage2[87]), .outData_88(wire_switch_out_stage2[88]), .outData_89(wire_switch_out_stage2[89]), .outData_90(wire_switch_out_stage2[90]), .outData_91(wire_switch_out_stage2[91]), .outData_92(wire_switch_out_stage2[92]), .outData_93(wire_switch_out_stage2[93]), .outData_94(wire_switch_out_stage2[94]), .outData_95(wire_switch_out_stage2[95]), .outData_96(wire_switch_out_stage2[96]), .outData_97(wire_switch_out_stage2[97]), .outData_98(wire_switch_out_stage2[98]), .outData_99(wire_switch_out_stage2[99]), .outData_100(wire_switch_out_stage2[100]), .outData_101(wire_switch_out_stage2[101]), .outData_102(wire_switch_out_stage2[102]), .outData_103(wire_switch_out_stage2[103]), .outData_104(wire_switch_out_stage2[104]), .outData_105(wire_switch_out_stage2[105]), .outData_106(wire_switch_out_stage2[106]), .outData_107(wire_switch_out_stage2[107]), .outData_108(wire_switch_out_stage2[108]), .outData_109(wire_switch_out_stage2[109]), .outData_110(wire_switch_out_stage2[110]), .outData_111(wire_switch_out_stage2[111]), .outData_112(wire_switch_out_stage2[112]), .outData_113(wire_switch_out_stage2[113]), .outData_114(wire_switch_out_stage2[114]), .outData_115(wire_switch_out_stage2[115]), .outData_116(wire_switch_out_stage2[116]), .outData_117(wire_switch_out_stage2[117]), .outData_118(wire_switch_out_stage2[118]), .outData_119(wire_switch_out_stage2[119]), .outData_120(wire_switch_out_stage2[120]), .outData_121(wire_switch_out_stage2[121]), .outData_122(wire_switch_out_stage2[122]), .outData_123(wire_switch_out_stage2[123]), .outData_124(wire_switch_out_stage2[124]), .outData_125(wire_switch_out_stage2[125]), .outData_126(wire_switch_out_stage2[126]), .outData_127(wire_switch_out_stage2[127]), .outData_128(wire_switch_out_stage2[128]), .outData_129(wire_switch_out_stage2[129]), .outData_130(wire_switch_out_stage2[130]), .outData_131(wire_switch_out_stage2[131]), .outData_132(wire_switch_out_stage2[132]), .outData_133(wire_switch_out_stage2[133]), .outData_134(wire_switch_out_stage2[134]), .outData_135(wire_switch_out_stage2[135]), .outData_136(wire_switch_out_stage2[136]), .outData_137(wire_switch_out_stage2[137]), .outData_138(wire_switch_out_stage2[138]), .outData_139(wire_switch_out_stage2[139]), .outData_140(wire_switch_out_stage2[140]), .outData_141(wire_switch_out_stage2[141]), .outData_142(wire_switch_out_stage2[142]), .outData_143(wire_switch_out_stage2[143]), .outData_144(wire_switch_out_stage2[144]), .outData_145(wire_switch_out_stage2[145]), .outData_146(wire_switch_out_stage2[146]), .outData_147(wire_switch_out_stage2[147]), .outData_148(wire_switch_out_stage2[148]), .outData_149(wire_switch_out_stage2[149]), .outData_150(wire_switch_out_stage2[150]), .outData_151(wire_switch_out_stage2[151]), .outData_152(wire_switch_out_stage2[152]), .outData_153(wire_switch_out_stage2[153]), .outData_154(wire_switch_out_stage2[154]), .outData_155(wire_switch_out_stage2[155]), .outData_156(wire_switch_out_stage2[156]), .outData_157(wire_switch_out_stage2[157]), .outData_158(wire_switch_out_stage2[158]), .outData_159(wire_switch_out_stage2[159]), .outData_160(wire_switch_out_stage2[160]), .outData_161(wire_switch_out_stage2[161]), .outData_162(wire_switch_out_stage2[162]), .outData_163(wire_switch_out_stage2[163]), .outData_164(wire_switch_out_stage2[164]), .outData_165(wire_switch_out_stage2[165]), .outData_166(wire_switch_out_stage2[166]), .outData_167(wire_switch_out_stage2[167]), .outData_168(wire_switch_out_stage2[168]), .outData_169(wire_switch_out_stage2[169]), .outData_170(wire_switch_out_stage2[170]), .outData_171(wire_switch_out_stage2[171]), .outData_172(wire_switch_out_stage2[172]), .outData_173(wire_switch_out_stage2[173]), .outData_174(wire_switch_out_stage2[174]), .outData_175(wire_switch_out_stage2[175]), .outData_176(wire_switch_out_stage2[176]), .outData_177(wire_switch_out_stage2[177]), .outData_178(wire_switch_out_stage2[178]), .outData_179(wire_switch_out_stage2[179]), .outData_180(wire_switch_out_stage2[180]), .outData_181(wire_switch_out_stage2[181]), .outData_182(wire_switch_out_stage2[182]), .outData_183(wire_switch_out_stage2[183]), .outData_184(wire_switch_out_stage2[184]), .outData_185(wire_switch_out_stage2[185]), .outData_186(wire_switch_out_stage2[186]), .outData_187(wire_switch_out_stage2[187]), .outData_188(wire_switch_out_stage2[188]), .outData_189(wire_switch_out_stage2[189]), .outData_190(wire_switch_out_stage2[190]), .outData_191(wire_switch_out_stage2[191]), .outData_192(wire_switch_out_stage2[192]), .outData_193(wire_switch_out_stage2[193]), .outData_194(wire_switch_out_stage2[194]), .outData_195(wire_switch_out_stage2[195]), .outData_196(wire_switch_out_stage2[196]), .outData_197(wire_switch_out_stage2[197]), .outData_198(wire_switch_out_stage2[198]), .outData_199(wire_switch_out_stage2[199]), .outData_200(wire_switch_out_stage2[200]), .outData_201(wire_switch_out_stage2[201]), .outData_202(wire_switch_out_stage2[202]), .outData_203(wire_switch_out_stage2[203]), .outData_204(wire_switch_out_stage2[204]), .outData_205(wire_switch_out_stage2[205]), .outData_206(wire_switch_out_stage2[206]), .outData_207(wire_switch_out_stage2[207]), .outData_208(wire_switch_out_stage2[208]), .outData_209(wire_switch_out_stage2[209]), .outData_210(wire_switch_out_stage2[210]), .outData_211(wire_switch_out_stage2[211]), .outData_212(wire_switch_out_stage2[212]), .outData_213(wire_switch_out_stage2[213]), .outData_214(wire_switch_out_stage2[214]), .outData_215(wire_switch_out_stage2[215]), .outData_216(wire_switch_out_stage2[216]), .outData_217(wire_switch_out_stage2[217]), .outData_218(wire_switch_out_stage2[218]), .outData_219(wire_switch_out_stage2[219]), .outData_220(wire_switch_out_stage2[220]), .outData_221(wire_switch_out_stage2[221]), .outData_222(wire_switch_out_stage2[222]), .outData_223(wire_switch_out_stage2[223]), .outData_224(wire_switch_out_stage2[224]), .outData_225(wire_switch_out_stage2[225]), .outData_226(wire_switch_out_stage2[226]), .outData_227(wire_switch_out_stage2[227]), .outData_228(wire_switch_out_stage2[228]), .outData_229(wire_switch_out_stage2[229]), .outData_230(wire_switch_out_stage2[230]), .outData_231(wire_switch_out_stage2[231]), .outData_232(wire_switch_out_stage2[232]), .outData_233(wire_switch_out_stage2[233]), .outData_234(wire_switch_out_stage2[234]), .outData_235(wire_switch_out_stage2[235]), .outData_236(wire_switch_out_stage2[236]), .outData_237(wire_switch_out_stage2[237]), .outData_238(wire_switch_out_stage2[238]), .outData_239(wire_switch_out_stage2[239]), .outData_240(wire_switch_out_stage2[240]), .outData_241(wire_switch_out_stage2[241]), .outData_242(wire_switch_out_stage2[242]), .outData_243(wire_switch_out_stage2[243]), .outData_244(wire_switch_out_stage2[244]), .outData_245(wire_switch_out_stage2[245]), .outData_246(wire_switch_out_stage2[246]), .outData_247(wire_switch_out_stage2[247]), .outData_248(wire_switch_out_stage2[248]), .outData_249(wire_switch_out_stage2[249]), .outData_250(wire_switch_out_stage2[250]), .outData_251(wire_switch_out_stage2[251]), .outData_252(wire_switch_out_stage2[252]), .outData_253(wire_switch_out_stage2[253]), .outData_254(wire_switch_out_stage2[254]), .outData_255(wire_switch_out_stage2[255]), 
        .in_start(con_in_start_stage2), .out_start(in_start_stage1), .ctrl(wire_ctrl_stage2), .clk(clk), .rst(rst));
  
  wireCon_dp256_st2_R wire_stage_2(
        .inData_0(wire_switch_out_stage3[0]), .inData_1(wire_switch_out_stage3[1]), .inData_2(wire_switch_out_stage3[2]), .inData_3(wire_switch_out_stage3[3]), .inData_4(wire_switch_out_stage3[4]), .inData_5(wire_switch_out_stage3[5]), .inData_6(wire_switch_out_stage3[6]), .inData_7(wire_switch_out_stage3[7]), .inData_8(wire_switch_out_stage3[8]), .inData_9(wire_switch_out_stage3[9]), .inData_10(wire_switch_out_stage3[10]), .inData_11(wire_switch_out_stage3[11]), .inData_12(wire_switch_out_stage3[12]), .inData_13(wire_switch_out_stage3[13]), .inData_14(wire_switch_out_stage3[14]), .inData_15(wire_switch_out_stage3[15]), .inData_16(wire_switch_out_stage3[16]), .inData_17(wire_switch_out_stage3[17]), .inData_18(wire_switch_out_stage3[18]), .inData_19(wire_switch_out_stage3[19]), .inData_20(wire_switch_out_stage3[20]), .inData_21(wire_switch_out_stage3[21]), .inData_22(wire_switch_out_stage3[22]), .inData_23(wire_switch_out_stage3[23]), .inData_24(wire_switch_out_stage3[24]), .inData_25(wire_switch_out_stage3[25]), .inData_26(wire_switch_out_stage3[26]), .inData_27(wire_switch_out_stage3[27]), .inData_28(wire_switch_out_stage3[28]), .inData_29(wire_switch_out_stage3[29]), .inData_30(wire_switch_out_stage3[30]), .inData_31(wire_switch_out_stage3[31]), .inData_32(wire_switch_out_stage3[32]), .inData_33(wire_switch_out_stage3[33]), .inData_34(wire_switch_out_stage3[34]), .inData_35(wire_switch_out_stage3[35]), .inData_36(wire_switch_out_stage3[36]), .inData_37(wire_switch_out_stage3[37]), .inData_38(wire_switch_out_stage3[38]), .inData_39(wire_switch_out_stage3[39]), .inData_40(wire_switch_out_stage3[40]), .inData_41(wire_switch_out_stage3[41]), .inData_42(wire_switch_out_stage3[42]), .inData_43(wire_switch_out_stage3[43]), .inData_44(wire_switch_out_stage3[44]), .inData_45(wire_switch_out_stage3[45]), .inData_46(wire_switch_out_stage3[46]), .inData_47(wire_switch_out_stage3[47]), .inData_48(wire_switch_out_stage3[48]), .inData_49(wire_switch_out_stage3[49]), .inData_50(wire_switch_out_stage3[50]), .inData_51(wire_switch_out_stage3[51]), .inData_52(wire_switch_out_stage3[52]), .inData_53(wire_switch_out_stage3[53]), .inData_54(wire_switch_out_stage3[54]), .inData_55(wire_switch_out_stage3[55]), .inData_56(wire_switch_out_stage3[56]), .inData_57(wire_switch_out_stage3[57]), .inData_58(wire_switch_out_stage3[58]), .inData_59(wire_switch_out_stage3[59]), .inData_60(wire_switch_out_stage3[60]), .inData_61(wire_switch_out_stage3[61]), .inData_62(wire_switch_out_stage3[62]), .inData_63(wire_switch_out_stage3[63]), .inData_64(wire_switch_out_stage3[64]), .inData_65(wire_switch_out_stage3[65]), .inData_66(wire_switch_out_stage3[66]), .inData_67(wire_switch_out_stage3[67]), .inData_68(wire_switch_out_stage3[68]), .inData_69(wire_switch_out_stage3[69]), .inData_70(wire_switch_out_stage3[70]), .inData_71(wire_switch_out_stage3[71]), .inData_72(wire_switch_out_stage3[72]), .inData_73(wire_switch_out_stage3[73]), .inData_74(wire_switch_out_stage3[74]), .inData_75(wire_switch_out_stage3[75]), .inData_76(wire_switch_out_stage3[76]), .inData_77(wire_switch_out_stage3[77]), .inData_78(wire_switch_out_stage3[78]), .inData_79(wire_switch_out_stage3[79]), .inData_80(wire_switch_out_stage3[80]), .inData_81(wire_switch_out_stage3[81]), .inData_82(wire_switch_out_stage3[82]), .inData_83(wire_switch_out_stage3[83]), .inData_84(wire_switch_out_stage3[84]), .inData_85(wire_switch_out_stage3[85]), .inData_86(wire_switch_out_stage3[86]), .inData_87(wire_switch_out_stage3[87]), .inData_88(wire_switch_out_stage3[88]), .inData_89(wire_switch_out_stage3[89]), .inData_90(wire_switch_out_stage3[90]), .inData_91(wire_switch_out_stage3[91]), .inData_92(wire_switch_out_stage3[92]), .inData_93(wire_switch_out_stage3[93]), .inData_94(wire_switch_out_stage3[94]), .inData_95(wire_switch_out_stage3[95]), .inData_96(wire_switch_out_stage3[96]), .inData_97(wire_switch_out_stage3[97]), .inData_98(wire_switch_out_stage3[98]), .inData_99(wire_switch_out_stage3[99]), .inData_100(wire_switch_out_stage3[100]), .inData_101(wire_switch_out_stage3[101]), .inData_102(wire_switch_out_stage3[102]), .inData_103(wire_switch_out_stage3[103]), .inData_104(wire_switch_out_stage3[104]), .inData_105(wire_switch_out_stage3[105]), .inData_106(wire_switch_out_stage3[106]), .inData_107(wire_switch_out_stage3[107]), .inData_108(wire_switch_out_stage3[108]), .inData_109(wire_switch_out_stage3[109]), .inData_110(wire_switch_out_stage3[110]), .inData_111(wire_switch_out_stage3[111]), .inData_112(wire_switch_out_stage3[112]), .inData_113(wire_switch_out_stage3[113]), .inData_114(wire_switch_out_stage3[114]), .inData_115(wire_switch_out_stage3[115]), .inData_116(wire_switch_out_stage3[116]), .inData_117(wire_switch_out_stage3[117]), .inData_118(wire_switch_out_stage3[118]), .inData_119(wire_switch_out_stage3[119]), .inData_120(wire_switch_out_stage3[120]), .inData_121(wire_switch_out_stage3[121]), .inData_122(wire_switch_out_stage3[122]), .inData_123(wire_switch_out_stage3[123]), .inData_124(wire_switch_out_stage3[124]), .inData_125(wire_switch_out_stage3[125]), .inData_126(wire_switch_out_stage3[126]), .inData_127(wire_switch_out_stage3[127]), .inData_128(wire_switch_out_stage3[128]), .inData_129(wire_switch_out_stage3[129]), .inData_130(wire_switch_out_stage3[130]), .inData_131(wire_switch_out_stage3[131]), .inData_132(wire_switch_out_stage3[132]), .inData_133(wire_switch_out_stage3[133]), .inData_134(wire_switch_out_stage3[134]), .inData_135(wire_switch_out_stage3[135]), .inData_136(wire_switch_out_stage3[136]), .inData_137(wire_switch_out_stage3[137]), .inData_138(wire_switch_out_stage3[138]), .inData_139(wire_switch_out_stage3[139]), .inData_140(wire_switch_out_stage3[140]), .inData_141(wire_switch_out_stage3[141]), .inData_142(wire_switch_out_stage3[142]), .inData_143(wire_switch_out_stage3[143]), .inData_144(wire_switch_out_stage3[144]), .inData_145(wire_switch_out_stage3[145]), .inData_146(wire_switch_out_stage3[146]), .inData_147(wire_switch_out_stage3[147]), .inData_148(wire_switch_out_stage3[148]), .inData_149(wire_switch_out_stage3[149]), .inData_150(wire_switch_out_stage3[150]), .inData_151(wire_switch_out_stage3[151]), .inData_152(wire_switch_out_stage3[152]), .inData_153(wire_switch_out_stage3[153]), .inData_154(wire_switch_out_stage3[154]), .inData_155(wire_switch_out_stage3[155]), .inData_156(wire_switch_out_stage3[156]), .inData_157(wire_switch_out_stage3[157]), .inData_158(wire_switch_out_stage3[158]), .inData_159(wire_switch_out_stage3[159]), .inData_160(wire_switch_out_stage3[160]), .inData_161(wire_switch_out_stage3[161]), .inData_162(wire_switch_out_stage3[162]), .inData_163(wire_switch_out_stage3[163]), .inData_164(wire_switch_out_stage3[164]), .inData_165(wire_switch_out_stage3[165]), .inData_166(wire_switch_out_stage3[166]), .inData_167(wire_switch_out_stage3[167]), .inData_168(wire_switch_out_stage3[168]), .inData_169(wire_switch_out_stage3[169]), .inData_170(wire_switch_out_stage3[170]), .inData_171(wire_switch_out_stage3[171]), .inData_172(wire_switch_out_stage3[172]), .inData_173(wire_switch_out_stage3[173]), .inData_174(wire_switch_out_stage3[174]), .inData_175(wire_switch_out_stage3[175]), .inData_176(wire_switch_out_stage3[176]), .inData_177(wire_switch_out_stage3[177]), .inData_178(wire_switch_out_stage3[178]), .inData_179(wire_switch_out_stage3[179]), .inData_180(wire_switch_out_stage3[180]), .inData_181(wire_switch_out_stage3[181]), .inData_182(wire_switch_out_stage3[182]), .inData_183(wire_switch_out_stage3[183]), .inData_184(wire_switch_out_stage3[184]), .inData_185(wire_switch_out_stage3[185]), .inData_186(wire_switch_out_stage3[186]), .inData_187(wire_switch_out_stage3[187]), .inData_188(wire_switch_out_stage3[188]), .inData_189(wire_switch_out_stage3[189]), .inData_190(wire_switch_out_stage3[190]), .inData_191(wire_switch_out_stage3[191]), .inData_192(wire_switch_out_stage3[192]), .inData_193(wire_switch_out_stage3[193]), .inData_194(wire_switch_out_stage3[194]), .inData_195(wire_switch_out_stage3[195]), .inData_196(wire_switch_out_stage3[196]), .inData_197(wire_switch_out_stage3[197]), .inData_198(wire_switch_out_stage3[198]), .inData_199(wire_switch_out_stage3[199]), .inData_200(wire_switch_out_stage3[200]), .inData_201(wire_switch_out_stage3[201]), .inData_202(wire_switch_out_stage3[202]), .inData_203(wire_switch_out_stage3[203]), .inData_204(wire_switch_out_stage3[204]), .inData_205(wire_switch_out_stage3[205]), .inData_206(wire_switch_out_stage3[206]), .inData_207(wire_switch_out_stage3[207]), .inData_208(wire_switch_out_stage3[208]), .inData_209(wire_switch_out_stage3[209]), .inData_210(wire_switch_out_stage3[210]), .inData_211(wire_switch_out_stage3[211]), .inData_212(wire_switch_out_stage3[212]), .inData_213(wire_switch_out_stage3[213]), .inData_214(wire_switch_out_stage3[214]), .inData_215(wire_switch_out_stage3[215]), .inData_216(wire_switch_out_stage3[216]), .inData_217(wire_switch_out_stage3[217]), .inData_218(wire_switch_out_stage3[218]), .inData_219(wire_switch_out_stage3[219]), .inData_220(wire_switch_out_stage3[220]), .inData_221(wire_switch_out_stage3[221]), .inData_222(wire_switch_out_stage3[222]), .inData_223(wire_switch_out_stage3[223]), .inData_224(wire_switch_out_stage3[224]), .inData_225(wire_switch_out_stage3[225]), .inData_226(wire_switch_out_stage3[226]), .inData_227(wire_switch_out_stage3[227]), .inData_228(wire_switch_out_stage3[228]), .inData_229(wire_switch_out_stage3[229]), .inData_230(wire_switch_out_stage3[230]), .inData_231(wire_switch_out_stage3[231]), .inData_232(wire_switch_out_stage3[232]), .inData_233(wire_switch_out_stage3[233]), .inData_234(wire_switch_out_stage3[234]), .inData_235(wire_switch_out_stage3[235]), .inData_236(wire_switch_out_stage3[236]), .inData_237(wire_switch_out_stage3[237]), .inData_238(wire_switch_out_stage3[238]), .inData_239(wire_switch_out_stage3[239]), .inData_240(wire_switch_out_stage3[240]), .inData_241(wire_switch_out_stage3[241]), .inData_242(wire_switch_out_stage3[242]), .inData_243(wire_switch_out_stage3[243]), .inData_244(wire_switch_out_stage3[244]), .inData_245(wire_switch_out_stage3[245]), .inData_246(wire_switch_out_stage3[246]), .inData_247(wire_switch_out_stage3[247]), .inData_248(wire_switch_out_stage3[248]), .inData_249(wire_switch_out_stage3[249]), .inData_250(wire_switch_out_stage3[250]), .inData_251(wire_switch_out_stage3[251]), .inData_252(wire_switch_out_stage3[252]), .inData_253(wire_switch_out_stage3[253]), .inData_254(wire_switch_out_stage3[254]), .inData_255(wire_switch_out_stage3[255]), 
        .outData_0(wire_switch_in_stage2[0]), .outData_1(wire_switch_in_stage2[1]), .outData_2(wire_switch_in_stage2[2]), .outData_3(wire_switch_in_stage2[3]), .outData_4(wire_switch_in_stage2[4]), .outData_5(wire_switch_in_stage2[5]), .outData_6(wire_switch_in_stage2[6]), .outData_7(wire_switch_in_stage2[7]), .outData_8(wire_switch_in_stage2[8]), .outData_9(wire_switch_in_stage2[9]), .outData_10(wire_switch_in_stage2[10]), .outData_11(wire_switch_in_stage2[11]), .outData_12(wire_switch_in_stage2[12]), .outData_13(wire_switch_in_stage2[13]), .outData_14(wire_switch_in_stage2[14]), .outData_15(wire_switch_in_stage2[15]), .outData_16(wire_switch_in_stage2[16]), .outData_17(wire_switch_in_stage2[17]), .outData_18(wire_switch_in_stage2[18]), .outData_19(wire_switch_in_stage2[19]), .outData_20(wire_switch_in_stage2[20]), .outData_21(wire_switch_in_stage2[21]), .outData_22(wire_switch_in_stage2[22]), .outData_23(wire_switch_in_stage2[23]), .outData_24(wire_switch_in_stage2[24]), .outData_25(wire_switch_in_stage2[25]), .outData_26(wire_switch_in_stage2[26]), .outData_27(wire_switch_in_stage2[27]), .outData_28(wire_switch_in_stage2[28]), .outData_29(wire_switch_in_stage2[29]), .outData_30(wire_switch_in_stage2[30]), .outData_31(wire_switch_in_stage2[31]), .outData_32(wire_switch_in_stage2[32]), .outData_33(wire_switch_in_stage2[33]), .outData_34(wire_switch_in_stage2[34]), .outData_35(wire_switch_in_stage2[35]), .outData_36(wire_switch_in_stage2[36]), .outData_37(wire_switch_in_stage2[37]), .outData_38(wire_switch_in_stage2[38]), .outData_39(wire_switch_in_stage2[39]), .outData_40(wire_switch_in_stage2[40]), .outData_41(wire_switch_in_stage2[41]), .outData_42(wire_switch_in_stage2[42]), .outData_43(wire_switch_in_stage2[43]), .outData_44(wire_switch_in_stage2[44]), .outData_45(wire_switch_in_stage2[45]), .outData_46(wire_switch_in_stage2[46]), .outData_47(wire_switch_in_stage2[47]), .outData_48(wire_switch_in_stage2[48]), .outData_49(wire_switch_in_stage2[49]), .outData_50(wire_switch_in_stage2[50]), .outData_51(wire_switch_in_stage2[51]), .outData_52(wire_switch_in_stage2[52]), .outData_53(wire_switch_in_stage2[53]), .outData_54(wire_switch_in_stage2[54]), .outData_55(wire_switch_in_stage2[55]), .outData_56(wire_switch_in_stage2[56]), .outData_57(wire_switch_in_stage2[57]), .outData_58(wire_switch_in_stage2[58]), .outData_59(wire_switch_in_stage2[59]), .outData_60(wire_switch_in_stage2[60]), .outData_61(wire_switch_in_stage2[61]), .outData_62(wire_switch_in_stage2[62]), .outData_63(wire_switch_in_stage2[63]), .outData_64(wire_switch_in_stage2[64]), .outData_65(wire_switch_in_stage2[65]), .outData_66(wire_switch_in_stage2[66]), .outData_67(wire_switch_in_stage2[67]), .outData_68(wire_switch_in_stage2[68]), .outData_69(wire_switch_in_stage2[69]), .outData_70(wire_switch_in_stage2[70]), .outData_71(wire_switch_in_stage2[71]), .outData_72(wire_switch_in_stage2[72]), .outData_73(wire_switch_in_stage2[73]), .outData_74(wire_switch_in_stage2[74]), .outData_75(wire_switch_in_stage2[75]), .outData_76(wire_switch_in_stage2[76]), .outData_77(wire_switch_in_stage2[77]), .outData_78(wire_switch_in_stage2[78]), .outData_79(wire_switch_in_stage2[79]), .outData_80(wire_switch_in_stage2[80]), .outData_81(wire_switch_in_stage2[81]), .outData_82(wire_switch_in_stage2[82]), .outData_83(wire_switch_in_stage2[83]), .outData_84(wire_switch_in_stage2[84]), .outData_85(wire_switch_in_stage2[85]), .outData_86(wire_switch_in_stage2[86]), .outData_87(wire_switch_in_stage2[87]), .outData_88(wire_switch_in_stage2[88]), .outData_89(wire_switch_in_stage2[89]), .outData_90(wire_switch_in_stage2[90]), .outData_91(wire_switch_in_stage2[91]), .outData_92(wire_switch_in_stage2[92]), .outData_93(wire_switch_in_stage2[93]), .outData_94(wire_switch_in_stage2[94]), .outData_95(wire_switch_in_stage2[95]), .outData_96(wire_switch_in_stage2[96]), .outData_97(wire_switch_in_stage2[97]), .outData_98(wire_switch_in_stage2[98]), .outData_99(wire_switch_in_stage2[99]), .outData_100(wire_switch_in_stage2[100]), .outData_101(wire_switch_in_stage2[101]), .outData_102(wire_switch_in_stage2[102]), .outData_103(wire_switch_in_stage2[103]), .outData_104(wire_switch_in_stage2[104]), .outData_105(wire_switch_in_stage2[105]), .outData_106(wire_switch_in_stage2[106]), .outData_107(wire_switch_in_stage2[107]), .outData_108(wire_switch_in_stage2[108]), .outData_109(wire_switch_in_stage2[109]), .outData_110(wire_switch_in_stage2[110]), .outData_111(wire_switch_in_stage2[111]), .outData_112(wire_switch_in_stage2[112]), .outData_113(wire_switch_in_stage2[113]), .outData_114(wire_switch_in_stage2[114]), .outData_115(wire_switch_in_stage2[115]), .outData_116(wire_switch_in_stage2[116]), .outData_117(wire_switch_in_stage2[117]), .outData_118(wire_switch_in_stage2[118]), .outData_119(wire_switch_in_stage2[119]), .outData_120(wire_switch_in_stage2[120]), .outData_121(wire_switch_in_stage2[121]), .outData_122(wire_switch_in_stage2[122]), .outData_123(wire_switch_in_stage2[123]), .outData_124(wire_switch_in_stage2[124]), .outData_125(wire_switch_in_stage2[125]), .outData_126(wire_switch_in_stage2[126]), .outData_127(wire_switch_in_stage2[127]), .outData_128(wire_switch_in_stage2[128]), .outData_129(wire_switch_in_stage2[129]), .outData_130(wire_switch_in_stage2[130]), .outData_131(wire_switch_in_stage2[131]), .outData_132(wire_switch_in_stage2[132]), .outData_133(wire_switch_in_stage2[133]), .outData_134(wire_switch_in_stage2[134]), .outData_135(wire_switch_in_stage2[135]), .outData_136(wire_switch_in_stage2[136]), .outData_137(wire_switch_in_stage2[137]), .outData_138(wire_switch_in_stage2[138]), .outData_139(wire_switch_in_stage2[139]), .outData_140(wire_switch_in_stage2[140]), .outData_141(wire_switch_in_stage2[141]), .outData_142(wire_switch_in_stage2[142]), .outData_143(wire_switch_in_stage2[143]), .outData_144(wire_switch_in_stage2[144]), .outData_145(wire_switch_in_stage2[145]), .outData_146(wire_switch_in_stage2[146]), .outData_147(wire_switch_in_stage2[147]), .outData_148(wire_switch_in_stage2[148]), .outData_149(wire_switch_in_stage2[149]), .outData_150(wire_switch_in_stage2[150]), .outData_151(wire_switch_in_stage2[151]), .outData_152(wire_switch_in_stage2[152]), .outData_153(wire_switch_in_stage2[153]), .outData_154(wire_switch_in_stage2[154]), .outData_155(wire_switch_in_stage2[155]), .outData_156(wire_switch_in_stage2[156]), .outData_157(wire_switch_in_stage2[157]), .outData_158(wire_switch_in_stage2[158]), .outData_159(wire_switch_in_stage2[159]), .outData_160(wire_switch_in_stage2[160]), .outData_161(wire_switch_in_stage2[161]), .outData_162(wire_switch_in_stage2[162]), .outData_163(wire_switch_in_stage2[163]), .outData_164(wire_switch_in_stage2[164]), .outData_165(wire_switch_in_stage2[165]), .outData_166(wire_switch_in_stage2[166]), .outData_167(wire_switch_in_stage2[167]), .outData_168(wire_switch_in_stage2[168]), .outData_169(wire_switch_in_stage2[169]), .outData_170(wire_switch_in_stage2[170]), .outData_171(wire_switch_in_stage2[171]), .outData_172(wire_switch_in_stage2[172]), .outData_173(wire_switch_in_stage2[173]), .outData_174(wire_switch_in_stage2[174]), .outData_175(wire_switch_in_stage2[175]), .outData_176(wire_switch_in_stage2[176]), .outData_177(wire_switch_in_stage2[177]), .outData_178(wire_switch_in_stage2[178]), .outData_179(wire_switch_in_stage2[179]), .outData_180(wire_switch_in_stage2[180]), .outData_181(wire_switch_in_stage2[181]), .outData_182(wire_switch_in_stage2[182]), .outData_183(wire_switch_in_stage2[183]), .outData_184(wire_switch_in_stage2[184]), .outData_185(wire_switch_in_stage2[185]), .outData_186(wire_switch_in_stage2[186]), .outData_187(wire_switch_in_stage2[187]), .outData_188(wire_switch_in_stage2[188]), .outData_189(wire_switch_in_stage2[189]), .outData_190(wire_switch_in_stage2[190]), .outData_191(wire_switch_in_stage2[191]), .outData_192(wire_switch_in_stage2[192]), .outData_193(wire_switch_in_stage2[193]), .outData_194(wire_switch_in_stage2[194]), .outData_195(wire_switch_in_stage2[195]), .outData_196(wire_switch_in_stage2[196]), .outData_197(wire_switch_in_stage2[197]), .outData_198(wire_switch_in_stage2[198]), .outData_199(wire_switch_in_stage2[199]), .outData_200(wire_switch_in_stage2[200]), .outData_201(wire_switch_in_stage2[201]), .outData_202(wire_switch_in_stage2[202]), .outData_203(wire_switch_in_stage2[203]), .outData_204(wire_switch_in_stage2[204]), .outData_205(wire_switch_in_stage2[205]), .outData_206(wire_switch_in_stage2[206]), .outData_207(wire_switch_in_stage2[207]), .outData_208(wire_switch_in_stage2[208]), .outData_209(wire_switch_in_stage2[209]), .outData_210(wire_switch_in_stage2[210]), .outData_211(wire_switch_in_stage2[211]), .outData_212(wire_switch_in_stage2[212]), .outData_213(wire_switch_in_stage2[213]), .outData_214(wire_switch_in_stage2[214]), .outData_215(wire_switch_in_stage2[215]), .outData_216(wire_switch_in_stage2[216]), .outData_217(wire_switch_in_stage2[217]), .outData_218(wire_switch_in_stage2[218]), .outData_219(wire_switch_in_stage2[219]), .outData_220(wire_switch_in_stage2[220]), .outData_221(wire_switch_in_stage2[221]), .outData_222(wire_switch_in_stage2[222]), .outData_223(wire_switch_in_stage2[223]), .outData_224(wire_switch_in_stage2[224]), .outData_225(wire_switch_in_stage2[225]), .outData_226(wire_switch_in_stage2[226]), .outData_227(wire_switch_in_stage2[227]), .outData_228(wire_switch_in_stage2[228]), .outData_229(wire_switch_in_stage2[229]), .outData_230(wire_switch_in_stage2[230]), .outData_231(wire_switch_in_stage2[231]), .outData_232(wire_switch_in_stage2[232]), .outData_233(wire_switch_in_stage2[233]), .outData_234(wire_switch_in_stage2[234]), .outData_235(wire_switch_in_stage2[235]), .outData_236(wire_switch_in_stage2[236]), .outData_237(wire_switch_in_stage2[237]), .outData_238(wire_switch_in_stage2[238]), .outData_239(wire_switch_in_stage2[239]), .outData_240(wire_switch_in_stage2[240]), .outData_241(wire_switch_in_stage2[241]), .outData_242(wire_switch_in_stage2[242]), .outData_243(wire_switch_in_stage2[243]), .outData_244(wire_switch_in_stage2[244]), .outData_245(wire_switch_in_stage2[245]), .outData_246(wire_switch_in_stage2[246]), .outData_247(wire_switch_in_stage2[247]), .outData_248(wire_switch_in_stage2[248]), .outData_249(wire_switch_in_stage2[249]), .outData_250(wire_switch_in_stage2[250]), .outData_251(wire_switch_in_stage2[251]), .outData_252(wire_switch_in_stage2[252]), .outData_253(wire_switch_in_stage2[253]), .outData_254(wire_switch_in_stage2[254]), .outData_255(wire_switch_in_stage2[255]), 
        .in_start(in_start_stage2), .out_start(con_in_start_stage2), .clk(clk), .rst(rst)); 

  
  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[0] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[1] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[2] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[3] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[4] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[5] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[6] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[7] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[8] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[9] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[10] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[11] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[12] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[13] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[14] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[15] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[16] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[17] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[18] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[19] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[20] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[21] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[22] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[23] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[24] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[25] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[26] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[27] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[28] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[29] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[30] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[31] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[32] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[33] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[34] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[35] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[36] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[37] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[38] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[39] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[40] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[41] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[42] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[43] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[44] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[45] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[46] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[47] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[48] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[49] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[50] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[51] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[52] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[53] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[54] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[55] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[56] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[57] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[58] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[59] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[60] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[61] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[62] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[63] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[64] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[65] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[66] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[67] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[68] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[69] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[70] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[71] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[72] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[73] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[74] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[75] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[76] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[77] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[78] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[79] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[80] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[81] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[82] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[83] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[84] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[85] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[86] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[87] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[88] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[89] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[90] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[91] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[92] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[93] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[94] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[95] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[96] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[97] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[98] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[99] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[100] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[101] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[102] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[103] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[104] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[105] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[106] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[107] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[108] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[109] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[110] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[111] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[112] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[113] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[114] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[115] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[116] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[117] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[118] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[119] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[120] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[121] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[122] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[123] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[124] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[125] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[126] <= counter_w[5]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage2[127] <= counter_w[5]; 
  end                            

  wire [DATA_WIDTH-1:0] wire_switch_in_stage1[255:0];
  wire [DATA_WIDTH-1:0] wire_switch_out_stage1[255:0];
  reg [127:0] wire_ctrl_stage1;

  switches_stage_st1_0_R switch_stage_1(
        .inData_0(wire_switch_in_stage1[0]), .inData_1(wire_switch_in_stage1[1]), .inData_2(wire_switch_in_stage1[2]), .inData_3(wire_switch_in_stage1[3]), .inData_4(wire_switch_in_stage1[4]), .inData_5(wire_switch_in_stage1[5]), .inData_6(wire_switch_in_stage1[6]), .inData_7(wire_switch_in_stage1[7]), .inData_8(wire_switch_in_stage1[8]), .inData_9(wire_switch_in_stage1[9]), .inData_10(wire_switch_in_stage1[10]), .inData_11(wire_switch_in_stage1[11]), .inData_12(wire_switch_in_stage1[12]), .inData_13(wire_switch_in_stage1[13]), .inData_14(wire_switch_in_stage1[14]), .inData_15(wire_switch_in_stage1[15]), .inData_16(wire_switch_in_stage1[16]), .inData_17(wire_switch_in_stage1[17]), .inData_18(wire_switch_in_stage1[18]), .inData_19(wire_switch_in_stage1[19]), .inData_20(wire_switch_in_stage1[20]), .inData_21(wire_switch_in_stage1[21]), .inData_22(wire_switch_in_stage1[22]), .inData_23(wire_switch_in_stage1[23]), .inData_24(wire_switch_in_stage1[24]), .inData_25(wire_switch_in_stage1[25]), .inData_26(wire_switch_in_stage1[26]), .inData_27(wire_switch_in_stage1[27]), .inData_28(wire_switch_in_stage1[28]), .inData_29(wire_switch_in_stage1[29]), .inData_30(wire_switch_in_stage1[30]), .inData_31(wire_switch_in_stage1[31]), .inData_32(wire_switch_in_stage1[32]), .inData_33(wire_switch_in_stage1[33]), .inData_34(wire_switch_in_stage1[34]), .inData_35(wire_switch_in_stage1[35]), .inData_36(wire_switch_in_stage1[36]), .inData_37(wire_switch_in_stage1[37]), .inData_38(wire_switch_in_stage1[38]), .inData_39(wire_switch_in_stage1[39]), .inData_40(wire_switch_in_stage1[40]), .inData_41(wire_switch_in_stage1[41]), .inData_42(wire_switch_in_stage1[42]), .inData_43(wire_switch_in_stage1[43]), .inData_44(wire_switch_in_stage1[44]), .inData_45(wire_switch_in_stage1[45]), .inData_46(wire_switch_in_stage1[46]), .inData_47(wire_switch_in_stage1[47]), .inData_48(wire_switch_in_stage1[48]), .inData_49(wire_switch_in_stage1[49]), .inData_50(wire_switch_in_stage1[50]), .inData_51(wire_switch_in_stage1[51]), .inData_52(wire_switch_in_stage1[52]), .inData_53(wire_switch_in_stage1[53]), .inData_54(wire_switch_in_stage1[54]), .inData_55(wire_switch_in_stage1[55]), .inData_56(wire_switch_in_stage1[56]), .inData_57(wire_switch_in_stage1[57]), .inData_58(wire_switch_in_stage1[58]), .inData_59(wire_switch_in_stage1[59]), .inData_60(wire_switch_in_stage1[60]), .inData_61(wire_switch_in_stage1[61]), .inData_62(wire_switch_in_stage1[62]), .inData_63(wire_switch_in_stage1[63]), .inData_64(wire_switch_in_stage1[64]), .inData_65(wire_switch_in_stage1[65]), .inData_66(wire_switch_in_stage1[66]), .inData_67(wire_switch_in_stage1[67]), .inData_68(wire_switch_in_stage1[68]), .inData_69(wire_switch_in_stage1[69]), .inData_70(wire_switch_in_stage1[70]), .inData_71(wire_switch_in_stage1[71]), .inData_72(wire_switch_in_stage1[72]), .inData_73(wire_switch_in_stage1[73]), .inData_74(wire_switch_in_stage1[74]), .inData_75(wire_switch_in_stage1[75]), .inData_76(wire_switch_in_stage1[76]), .inData_77(wire_switch_in_stage1[77]), .inData_78(wire_switch_in_stage1[78]), .inData_79(wire_switch_in_stage1[79]), .inData_80(wire_switch_in_stage1[80]), .inData_81(wire_switch_in_stage1[81]), .inData_82(wire_switch_in_stage1[82]), .inData_83(wire_switch_in_stage1[83]), .inData_84(wire_switch_in_stage1[84]), .inData_85(wire_switch_in_stage1[85]), .inData_86(wire_switch_in_stage1[86]), .inData_87(wire_switch_in_stage1[87]), .inData_88(wire_switch_in_stage1[88]), .inData_89(wire_switch_in_stage1[89]), .inData_90(wire_switch_in_stage1[90]), .inData_91(wire_switch_in_stage1[91]), .inData_92(wire_switch_in_stage1[92]), .inData_93(wire_switch_in_stage1[93]), .inData_94(wire_switch_in_stage1[94]), .inData_95(wire_switch_in_stage1[95]), .inData_96(wire_switch_in_stage1[96]), .inData_97(wire_switch_in_stage1[97]), .inData_98(wire_switch_in_stage1[98]), .inData_99(wire_switch_in_stage1[99]), .inData_100(wire_switch_in_stage1[100]), .inData_101(wire_switch_in_stage1[101]), .inData_102(wire_switch_in_stage1[102]), .inData_103(wire_switch_in_stage1[103]), .inData_104(wire_switch_in_stage1[104]), .inData_105(wire_switch_in_stage1[105]), .inData_106(wire_switch_in_stage1[106]), .inData_107(wire_switch_in_stage1[107]), .inData_108(wire_switch_in_stage1[108]), .inData_109(wire_switch_in_stage1[109]), .inData_110(wire_switch_in_stage1[110]), .inData_111(wire_switch_in_stage1[111]), .inData_112(wire_switch_in_stage1[112]), .inData_113(wire_switch_in_stage1[113]), .inData_114(wire_switch_in_stage1[114]), .inData_115(wire_switch_in_stage1[115]), .inData_116(wire_switch_in_stage1[116]), .inData_117(wire_switch_in_stage1[117]), .inData_118(wire_switch_in_stage1[118]), .inData_119(wire_switch_in_stage1[119]), .inData_120(wire_switch_in_stage1[120]), .inData_121(wire_switch_in_stage1[121]), .inData_122(wire_switch_in_stage1[122]), .inData_123(wire_switch_in_stage1[123]), .inData_124(wire_switch_in_stage1[124]), .inData_125(wire_switch_in_stage1[125]), .inData_126(wire_switch_in_stage1[126]), .inData_127(wire_switch_in_stage1[127]), .inData_128(wire_switch_in_stage1[128]), .inData_129(wire_switch_in_stage1[129]), .inData_130(wire_switch_in_stage1[130]), .inData_131(wire_switch_in_stage1[131]), .inData_132(wire_switch_in_stage1[132]), .inData_133(wire_switch_in_stage1[133]), .inData_134(wire_switch_in_stage1[134]), .inData_135(wire_switch_in_stage1[135]), .inData_136(wire_switch_in_stage1[136]), .inData_137(wire_switch_in_stage1[137]), .inData_138(wire_switch_in_stage1[138]), .inData_139(wire_switch_in_stage1[139]), .inData_140(wire_switch_in_stage1[140]), .inData_141(wire_switch_in_stage1[141]), .inData_142(wire_switch_in_stage1[142]), .inData_143(wire_switch_in_stage1[143]), .inData_144(wire_switch_in_stage1[144]), .inData_145(wire_switch_in_stage1[145]), .inData_146(wire_switch_in_stage1[146]), .inData_147(wire_switch_in_stage1[147]), .inData_148(wire_switch_in_stage1[148]), .inData_149(wire_switch_in_stage1[149]), .inData_150(wire_switch_in_stage1[150]), .inData_151(wire_switch_in_stage1[151]), .inData_152(wire_switch_in_stage1[152]), .inData_153(wire_switch_in_stage1[153]), .inData_154(wire_switch_in_stage1[154]), .inData_155(wire_switch_in_stage1[155]), .inData_156(wire_switch_in_stage1[156]), .inData_157(wire_switch_in_stage1[157]), .inData_158(wire_switch_in_stage1[158]), .inData_159(wire_switch_in_stage1[159]), .inData_160(wire_switch_in_stage1[160]), .inData_161(wire_switch_in_stage1[161]), .inData_162(wire_switch_in_stage1[162]), .inData_163(wire_switch_in_stage1[163]), .inData_164(wire_switch_in_stage1[164]), .inData_165(wire_switch_in_stage1[165]), .inData_166(wire_switch_in_stage1[166]), .inData_167(wire_switch_in_stage1[167]), .inData_168(wire_switch_in_stage1[168]), .inData_169(wire_switch_in_stage1[169]), .inData_170(wire_switch_in_stage1[170]), .inData_171(wire_switch_in_stage1[171]), .inData_172(wire_switch_in_stage1[172]), .inData_173(wire_switch_in_stage1[173]), .inData_174(wire_switch_in_stage1[174]), .inData_175(wire_switch_in_stage1[175]), .inData_176(wire_switch_in_stage1[176]), .inData_177(wire_switch_in_stage1[177]), .inData_178(wire_switch_in_stage1[178]), .inData_179(wire_switch_in_stage1[179]), .inData_180(wire_switch_in_stage1[180]), .inData_181(wire_switch_in_stage1[181]), .inData_182(wire_switch_in_stage1[182]), .inData_183(wire_switch_in_stage1[183]), .inData_184(wire_switch_in_stage1[184]), .inData_185(wire_switch_in_stage1[185]), .inData_186(wire_switch_in_stage1[186]), .inData_187(wire_switch_in_stage1[187]), .inData_188(wire_switch_in_stage1[188]), .inData_189(wire_switch_in_stage1[189]), .inData_190(wire_switch_in_stage1[190]), .inData_191(wire_switch_in_stage1[191]), .inData_192(wire_switch_in_stage1[192]), .inData_193(wire_switch_in_stage1[193]), .inData_194(wire_switch_in_stage1[194]), .inData_195(wire_switch_in_stage1[195]), .inData_196(wire_switch_in_stage1[196]), .inData_197(wire_switch_in_stage1[197]), .inData_198(wire_switch_in_stage1[198]), .inData_199(wire_switch_in_stage1[199]), .inData_200(wire_switch_in_stage1[200]), .inData_201(wire_switch_in_stage1[201]), .inData_202(wire_switch_in_stage1[202]), .inData_203(wire_switch_in_stage1[203]), .inData_204(wire_switch_in_stage1[204]), .inData_205(wire_switch_in_stage1[205]), .inData_206(wire_switch_in_stage1[206]), .inData_207(wire_switch_in_stage1[207]), .inData_208(wire_switch_in_stage1[208]), .inData_209(wire_switch_in_stage1[209]), .inData_210(wire_switch_in_stage1[210]), .inData_211(wire_switch_in_stage1[211]), .inData_212(wire_switch_in_stage1[212]), .inData_213(wire_switch_in_stage1[213]), .inData_214(wire_switch_in_stage1[214]), .inData_215(wire_switch_in_stage1[215]), .inData_216(wire_switch_in_stage1[216]), .inData_217(wire_switch_in_stage1[217]), .inData_218(wire_switch_in_stage1[218]), .inData_219(wire_switch_in_stage1[219]), .inData_220(wire_switch_in_stage1[220]), .inData_221(wire_switch_in_stage1[221]), .inData_222(wire_switch_in_stage1[222]), .inData_223(wire_switch_in_stage1[223]), .inData_224(wire_switch_in_stage1[224]), .inData_225(wire_switch_in_stage1[225]), .inData_226(wire_switch_in_stage1[226]), .inData_227(wire_switch_in_stage1[227]), .inData_228(wire_switch_in_stage1[228]), .inData_229(wire_switch_in_stage1[229]), .inData_230(wire_switch_in_stage1[230]), .inData_231(wire_switch_in_stage1[231]), .inData_232(wire_switch_in_stage1[232]), .inData_233(wire_switch_in_stage1[233]), .inData_234(wire_switch_in_stage1[234]), .inData_235(wire_switch_in_stage1[235]), .inData_236(wire_switch_in_stage1[236]), .inData_237(wire_switch_in_stage1[237]), .inData_238(wire_switch_in_stage1[238]), .inData_239(wire_switch_in_stage1[239]), .inData_240(wire_switch_in_stage1[240]), .inData_241(wire_switch_in_stage1[241]), .inData_242(wire_switch_in_stage1[242]), .inData_243(wire_switch_in_stage1[243]), .inData_244(wire_switch_in_stage1[244]), .inData_245(wire_switch_in_stage1[245]), .inData_246(wire_switch_in_stage1[246]), .inData_247(wire_switch_in_stage1[247]), .inData_248(wire_switch_in_stage1[248]), .inData_249(wire_switch_in_stage1[249]), .inData_250(wire_switch_in_stage1[250]), .inData_251(wire_switch_in_stage1[251]), .inData_252(wire_switch_in_stage1[252]), .inData_253(wire_switch_in_stage1[253]), .inData_254(wire_switch_in_stage1[254]), .inData_255(wire_switch_in_stage1[255]), 
        .outData_0(wire_switch_out_stage1[0]), .outData_1(wire_switch_out_stage1[1]), .outData_2(wire_switch_out_stage1[2]), .outData_3(wire_switch_out_stage1[3]), .outData_4(wire_switch_out_stage1[4]), .outData_5(wire_switch_out_stage1[5]), .outData_6(wire_switch_out_stage1[6]), .outData_7(wire_switch_out_stage1[7]), .outData_8(wire_switch_out_stage1[8]), .outData_9(wire_switch_out_stage1[9]), .outData_10(wire_switch_out_stage1[10]), .outData_11(wire_switch_out_stage1[11]), .outData_12(wire_switch_out_stage1[12]), .outData_13(wire_switch_out_stage1[13]), .outData_14(wire_switch_out_stage1[14]), .outData_15(wire_switch_out_stage1[15]), .outData_16(wire_switch_out_stage1[16]), .outData_17(wire_switch_out_stage1[17]), .outData_18(wire_switch_out_stage1[18]), .outData_19(wire_switch_out_stage1[19]), .outData_20(wire_switch_out_stage1[20]), .outData_21(wire_switch_out_stage1[21]), .outData_22(wire_switch_out_stage1[22]), .outData_23(wire_switch_out_stage1[23]), .outData_24(wire_switch_out_stage1[24]), .outData_25(wire_switch_out_stage1[25]), .outData_26(wire_switch_out_stage1[26]), .outData_27(wire_switch_out_stage1[27]), .outData_28(wire_switch_out_stage1[28]), .outData_29(wire_switch_out_stage1[29]), .outData_30(wire_switch_out_stage1[30]), .outData_31(wire_switch_out_stage1[31]), .outData_32(wire_switch_out_stage1[32]), .outData_33(wire_switch_out_stage1[33]), .outData_34(wire_switch_out_stage1[34]), .outData_35(wire_switch_out_stage1[35]), .outData_36(wire_switch_out_stage1[36]), .outData_37(wire_switch_out_stage1[37]), .outData_38(wire_switch_out_stage1[38]), .outData_39(wire_switch_out_stage1[39]), .outData_40(wire_switch_out_stage1[40]), .outData_41(wire_switch_out_stage1[41]), .outData_42(wire_switch_out_stage1[42]), .outData_43(wire_switch_out_stage1[43]), .outData_44(wire_switch_out_stage1[44]), .outData_45(wire_switch_out_stage1[45]), .outData_46(wire_switch_out_stage1[46]), .outData_47(wire_switch_out_stage1[47]), .outData_48(wire_switch_out_stage1[48]), .outData_49(wire_switch_out_stage1[49]), .outData_50(wire_switch_out_stage1[50]), .outData_51(wire_switch_out_stage1[51]), .outData_52(wire_switch_out_stage1[52]), .outData_53(wire_switch_out_stage1[53]), .outData_54(wire_switch_out_stage1[54]), .outData_55(wire_switch_out_stage1[55]), .outData_56(wire_switch_out_stage1[56]), .outData_57(wire_switch_out_stage1[57]), .outData_58(wire_switch_out_stage1[58]), .outData_59(wire_switch_out_stage1[59]), .outData_60(wire_switch_out_stage1[60]), .outData_61(wire_switch_out_stage1[61]), .outData_62(wire_switch_out_stage1[62]), .outData_63(wire_switch_out_stage1[63]), .outData_64(wire_switch_out_stage1[64]), .outData_65(wire_switch_out_stage1[65]), .outData_66(wire_switch_out_stage1[66]), .outData_67(wire_switch_out_stage1[67]), .outData_68(wire_switch_out_stage1[68]), .outData_69(wire_switch_out_stage1[69]), .outData_70(wire_switch_out_stage1[70]), .outData_71(wire_switch_out_stage1[71]), .outData_72(wire_switch_out_stage1[72]), .outData_73(wire_switch_out_stage1[73]), .outData_74(wire_switch_out_stage1[74]), .outData_75(wire_switch_out_stage1[75]), .outData_76(wire_switch_out_stage1[76]), .outData_77(wire_switch_out_stage1[77]), .outData_78(wire_switch_out_stage1[78]), .outData_79(wire_switch_out_stage1[79]), .outData_80(wire_switch_out_stage1[80]), .outData_81(wire_switch_out_stage1[81]), .outData_82(wire_switch_out_stage1[82]), .outData_83(wire_switch_out_stage1[83]), .outData_84(wire_switch_out_stage1[84]), .outData_85(wire_switch_out_stage1[85]), .outData_86(wire_switch_out_stage1[86]), .outData_87(wire_switch_out_stage1[87]), .outData_88(wire_switch_out_stage1[88]), .outData_89(wire_switch_out_stage1[89]), .outData_90(wire_switch_out_stage1[90]), .outData_91(wire_switch_out_stage1[91]), .outData_92(wire_switch_out_stage1[92]), .outData_93(wire_switch_out_stage1[93]), .outData_94(wire_switch_out_stage1[94]), .outData_95(wire_switch_out_stage1[95]), .outData_96(wire_switch_out_stage1[96]), .outData_97(wire_switch_out_stage1[97]), .outData_98(wire_switch_out_stage1[98]), .outData_99(wire_switch_out_stage1[99]), .outData_100(wire_switch_out_stage1[100]), .outData_101(wire_switch_out_stage1[101]), .outData_102(wire_switch_out_stage1[102]), .outData_103(wire_switch_out_stage1[103]), .outData_104(wire_switch_out_stage1[104]), .outData_105(wire_switch_out_stage1[105]), .outData_106(wire_switch_out_stage1[106]), .outData_107(wire_switch_out_stage1[107]), .outData_108(wire_switch_out_stage1[108]), .outData_109(wire_switch_out_stage1[109]), .outData_110(wire_switch_out_stage1[110]), .outData_111(wire_switch_out_stage1[111]), .outData_112(wire_switch_out_stage1[112]), .outData_113(wire_switch_out_stage1[113]), .outData_114(wire_switch_out_stage1[114]), .outData_115(wire_switch_out_stage1[115]), .outData_116(wire_switch_out_stage1[116]), .outData_117(wire_switch_out_stage1[117]), .outData_118(wire_switch_out_stage1[118]), .outData_119(wire_switch_out_stage1[119]), .outData_120(wire_switch_out_stage1[120]), .outData_121(wire_switch_out_stage1[121]), .outData_122(wire_switch_out_stage1[122]), .outData_123(wire_switch_out_stage1[123]), .outData_124(wire_switch_out_stage1[124]), .outData_125(wire_switch_out_stage1[125]), .outData_126(wire_switch_out_stage1[126]), .outData_127(wire_switch_out_stage1[127]), .outData_128(wire_switch_out_stage1[128]), .outData_129(wire_switch_out_stage1[129]), .outData_130(wire_switch_out_stage1[130]), .outData_131(wire_switch_out_stage1[131]), .outData_132(wire_switch_out_stage1[132]), .outData_133(wire_switch_out_stage1[133]), .outData_134(wire_switch_out_stage1[134]), .outData_135(wire_switch_out_stage1[135]), .outData_136(wire_switch_out_stage1[136]), .outData_137(wire_switch_out_stage1[137]), .outData_138(wire_switch_out_stage1[138]), .outData_139(wire_switch_out_stage1[139]), .outData_140(wire_switch_out_stage1[140]), .outData_141(wire_switch_out_stage1[141]), .outData_142(wire_switch_out_stage1[142]), .outData_143(wire_switch_out_stage1[143]), .outData_144(wire_switch_out_stage1[144]), .outData_145(wire_switch_out_stage1[145]), .outData_146(wire_switch_out_stage1[146]), .outData_147(wire_switch_out_stage1[147]), .outData_148(wire_switch_out_stage1[148]), .outData_149(wire_switch_out_stage1[149]), .outData_150(wire_switch_out_stage1[150]), .outData_151(wire_switch_out_stage1[151]), .outData_152(wire_switch_out_stage1[152]), .outData_153(wire_switch_out_stage1[153]), .outData_154(wire_switch_out_stage1[154]), .outData_155(wire_switch_out_stage1[155]), .outData_156(wire_switch_out_stage1[156]), .outData_157(wire_switch_out_stage1[157]), .outData_158(wire_switch_out_stage1[158]), .outData_159(wire_switch_out_stage1[159]), .outData_160(wire_switch_out_stage1[160]), .outData_161(wire_switch_out_stage1[161]), .outData_162(wire_switch_out_stage1[162]), .outData_163(wire_switch_out_stage1[163]), .outData_164(wire_switch_out_stage1[164]), .outData_165(wire_switch_out_stage1[165]), .outData_166(wire_switch_out_stage1[166]), .outData_167(wire_switch_out_stage1[167]), .outData_168(wire_switch_out_stage1[168]), .outData_169(wire_switch_out_stage1[169]), .outData_170(wire_switch_out_stage1[170]), .outData_171(wire_switch_out_stage1[171]), .outData_172(wire_switch_out_stage1[172]), .outData_173(wire_switch_out_stage1[173]), .outData_174(wire_switch_out_stage1[174]), .outData_175(wire_switch_out_stage1[175]), .outData_176(wire_switch_out_stage1[176]), .outData_177(wire_switch_out_stage1[177]), .outData_178(wire_switch_out_stage1[178]), .outData_179(wire_switch_out_stage1[179]), .outData_180(wire_switch_out_stage1[180]), .outData_181(wire_switch_out_stage1[181]), .outData_182(wire_switch_out_stage1[182]), .outData_183(wire_switch_out_stage1[183]), .outData_184(wire_switch_out_stage1[184]), .outData_185(wire_switch_out_stage1[185]), .outData_186(wire_switch_out_stage1[186]), .outData_187(wire_switch_out_stage1[187]), .outData_188(wire_switch_out_stage1[188]), .outData_189(wire_switch_out_stage1[189]), .outData_190(wire_switch_out_stage1[190]), .outData_191(wire_switch_out_stage1[191]), .outData_192(wire_switch_out_stage1[192]), .outData_193(wire_switch_out_stage1[193]), .outData_194(wire_switch_out_stage1[194]), .outData_195(wire_switch_out_stage1[195]), .outData_196(wire_switch_out_stage1[196]), .outData_197(wire_switch_out_stage1[197]), .outData_198(wire_switch_out_stage1[198]), .outData_199(wire_switch_out_stage1[199]), .outData_200(wire_switch_out_stage1[200]), .outData_201(wire_switch_out_stage1[201]), .outData_202(wire_switch_out_stage1[202]), .outData_203(wire_switch_out_stage1[203]), .outData_204(wire_switch_out_stage1[204]), .outData_205(wire_switch_out_stage1[205]), .outData_206(wire_switch_out_stage1[206]), .outData_207(wire_switch_out_stage1[207]), .outData_208(wire_switch_out_stage1[208]), .outData_209(wire_switch_out_stage1[209]), .outData_210(wire_switch_out_stage1[210]), .outData_211(wire_switch_out_stage1[211]), .outData_212(wire_switch_out_stage1[212]), .outData_213(wire_switch_out_stage1[213]), .outData_214(wire_switch_out_stage1[214]), .outData_215(wire_switch_out_stage1[215]), .outData_216(wire_switch_out_stage1[216]), .outData_217(wire_switch_out_stage1[217]), .outData_218(wire_switch_out_stage1[218]), .outData_219(wire_switch_out_stage1[219]), .outData_220(wire_switch_out_stage1[220]), .outData_221(wire_switch_out_stage1[221]), .outData_222(wire_switch_out_stage1[222]), .outData_223(wire_switch_out_stage1[223]), .outData_224(wire_switch_out_stage1[224]), .outData_225(wire_switch_out_stage1[225]), .outData_226(wire_switch_out_stage1[226]), .outData_227(wire_switch_out_stage1[227]), .outData_228(wire_switch_out_stage1[228]), .outData_229(wire_switch_out_stage1[229]), .outData_230(wire_switch_out_stage1[230]), .outData_231(wire_switch_out_stage1[231]), .outData_232(wire_switch_out_stage1[232]), .outData_233(wire_switch_out_stage1[233]), .outData_234(wire_switch_out_stage1[234]), .outData_235(wire_switch_out_stage1[235]), .outData_236(wire_switch_out_stage1[236]), .outData_237(wire_switch_out_stage1[237]), .outData_238(wire_switch_out_stage1[238]), .outData_239(wire_switch_out_stage1[239]), .outData_240(wire_switch_out_stage1[240]), .outData_241(wire_switch_out_stage1[241]), .outData_242(wire_switch_out_stage1[242]), .outData_243(wire_switch_out_stage1[243]), .outData_244(wire_switch_out_stage1[244]), .outData_245(wire_switch_out_stage1[245]), .outData_246(wire_switch_out_stage1[246]), .outData_247(wire_switch_out_stage1[247]), .outData_248(wire_switch_out_stage1[248]), .outData_249(wire_switch_out_stage1[249]), .outData_250(wire_switch_out_stage1[250]), .outData_251(wire_switch_out_stage1[251]), .outData_252(wire_switch_out_stage1[252]), .outData_253(wire_switch_out_stage1[253]), .outData_254(wire_switch_out_stage1[254]), .outData_255(wire_switch_out_stage1[255]), 
        .in_start(con_in_start_stage1), .out_start(in_start_stage0), .ctrl(wire_ctrl_stage1), .clk(clk), .rst(rst));
  
  wireCon_dp256_st1_R wire_stage_1(
        .inData_0(wire_switch_out_stage2[0]), .inData_1(wire_switch_out_stage2[1]), .inData_2(wire_switch_out_stage2[2]), .inData_3(wire_switch_out_stage2[3]), .inData_4(wire_switch_out_stage2[4]), .inData_5(wire_switch_out_stage2[5]), .inData_6(wire_switch_out_stage2[6]), .inData_7(wire_switch_out_stage2[7]), .inData_8(wire_switch_out_stage2[8]), .inData_9(wire_switch_out_stage2[9]), .inData_10(wire_switch_out_stage2[10]), .inData_11(wire_switch_out_stage2[11]), .inData_12(wire_switch_out_stage2[12]), .inData_13(wire_switch_out_stage2[13]), .inData_14(wire_switch_out_stage2[14]), .inData_15(wire_switch_out_stage2[15]), .inData_16(wire_switch_out_stage2[16]), .inData_17(wire_switch_out_stage2[17]), .inData_18(wire_switch_out_stage2[18]), .inData_19(wire_switch_out_stage2[19]), .inData_20(wire_switch_out_stage2[20]), .inData_21(wire_switch_out_stage2[21]), .inData_22(wire_switch_out_stage2[22]), .inData_23(wire_switch_out_stage2[23]), .inData_24(wire_switch_out_stage2[24]), .inData_25(wire_switch_out_stage2[25]), .inData_26(wire_switch_out_stage2[26]), .inData_27(wire_switch_out_stage2[27]), .inData_28(wire_switch_out_stage2[28]), .inData_29(wire_switch_out_stage2[29]), .inData_30(wire_switch_out_stage2[30]), .inData_31(wire_switch_out_stage2[31]), .inData_32(wire_switch_out_stage2[32]), .inData_33(wire_switch_out_stage2[33]), .inData_34(wire_switch_out_stage2[34]), .inData_35(wire_switch_out_stage2[35]), .inData_36(wire_switch_out_stage2[36]), .inData_37(wire_switch_out_stage2[37]), .inData_38(wire_switch_out_stage2[38]), .inData_39(wire_switch_out_stage2[39]), .inData_40(wire_switch_out_stage2[40]), .inData_41(wire_switch_out_stage2[41]), .inData_42(wire_switch_out_stage2[42]), .inData_43(wire_switch_out_stage2[43]), .inData_44(wire_switch_out_stage2[44]), .inData_45(wire_switch_out_stage2[45]), .inData_46(wire_switch_out_stage2[46]), .inData_47(wire_switch_out_stage2[47]), .inData_48(wire_switch_out_stage2[48]), .inData_49(wire_switch_out_stage2[49]), .inData_50(wire_switch_out_stage2[50]), .inData_51(wire_switch_out_stage2[51]), .inData_52(wire_switch_out_stage2[52]), .inData_53(wire_switch_out_stage2[53]), .inData_54(wire_switch_out_stage2[54]), .inData_55(wire_switch_out_stage2[55]), .inData_56(wire_switch_out_stage2[56]), .inData_57(wire_switch_out_stage2[57]), .inData_58(wire_switch_out_stage2[58]), .inData_59(wire_switch_out_stage2[59]), .inData_60(wire_switch_out_stage2[60]), .inData_61(wire_switch_out_stage2[61]), .inData_62(wire_switch_out_stage2[62]), .inData_63(wire_switch_out_stage2[63]), .inData_64(wire_switch_out_stage2[64]), .inData_65(wire_switch_out_stage2[65]), .inData_66(wire_switch_out_stage2[66]), .inData_67(wire_switch_out_stage2[67]), .inData_68(wire_switch_out_stage2[68]), .inData_69(wire_switch_out_stage2[69]), .inData_70(wire_switch_out_stage2[70]), .inData_71(wire_switch_out_stage2[71]), .inData_72(wire_switch_out_stage2[72]), .inData_73(wire_switch_out_stage2[73]), .inData_74(wire_switch_out_stage2[74]), .inData_75(wire_switch_out_stage2[75]), .inData_76(wire_switch_out_stage2[76]), .inData_77(wire_switch_out_stage2[77]), .inData_78(wire_switch_out_stage2[78]), .inData_79(wire_switch_out_stage2[79]), .inData_80(wire_switch_out_stage2[80]), .inData_81(wire_switch_out_stage2[81]), .inData_82(wire_switch_out_stage2[82]), .inData_83(wire_switch_out_stage2[83]), .inData_84(wire_switch_out_stage2[84]), .inData_85(wire_switch_out_stage2[85]), .inData_86(wire_switch_out_stage2[86]), .inData_87(wire_switch_out_stage2[87]), .inData_88(wire_switch_out_stage2[88]), .inData_89(wire_switch_out_stage2[89]), .inData_90(wire_switch_out_stage2[90]), .inData_91(wire_switch_out_stage2[91]), .inData_92(wire_switch_out_stage2[92]), .inData_93(wire_switch_out_stage2[93]), .inData_94(wire_switch_out_stage2[94]), .inData_95(wire_switch_out_stage2[95]), .inData_96(wire_switch_out_stage2[96]), .inData_97(wire_switch_out_stage2[97]), .inData_98(wire_switch_out_stage2[98]), .inData_99(wire_switch_out_stage2[99]), .inData_100(wire_switch_out_stage2[100]), .inData_101(wire_switch_out_stage2[101]), .inData_102(wire_switch_out_stage2[102]), .inData_103(wire_switch_out_stage2[103]), .inData_104(wire_switch_out_stage2[104]), .inData_105(wire_switch_out_stage2[105]), .inData_106(wire_switch_out_stage2[106]), .inData_107(wire_switch_out_stage2[107]), .inData_108(wire_switch_out_stage2[108]), .inData_109(wire_switch_out_stage2[109]), .inData_110(wire_switch_out_stage2[110]), .inData_111(wire_switch_out_stage2[111]), .inData_112(wire_switch_out_stage2[112]), .inData_113(wire_switch_out_stage2[113]), .inData_114(wire_switch_out_stage2[114]), .inData_115(wire_switch_out_stage2[115]), .inData_116(wire_switch_out_stage2[116]), .inData_117(wire_switch_out_stage2[117]), .inData_118(wire_switch_out_stage2[118]), .inData_119(wire_switch_out_stage2[119]), .inData_120(wire_switch_out_stage2[120]), .inData_121(wire_switch_out_stage2[121]), .inData_122(wire_switch_out_stage2[122]), .inData_123(wire_switch_out_stage2[123]), .inData_124(wire_switch_out_stage2[124]), .inData_125(wire_switch_out_stage2[125]), .inData_126(wire_switch_out_stage2[126]), .inData_127(wire_switch_out_stage2[127]), .inData_128(wire_switch_out_stage2[128]), .inData_129(wire_switch_out_stage2[129]), .inData_130(wire_switch_out_stage2[130]), .inData_131(wire_switch_out_stage2[131]), .inData_132(wire_switch_out_stage2[132]), .inData_133(wire_switch_out_stage2[133]), .inData_134(wire_switch_out_stage2[134]), .inData_135(wire_switch_out_stage2[135]), .inData_136(wire_switch_out_stage2[136]), .inData_137(wire_switch_out_stage2[137]), .inData_138(wire_switch_out_stage2[138]), .inData_139(wire_switch_out_stage2[139]), .inData_140(wire_switch_out_stage2[140]), .inData_141(wire_switch_out_stage2[141]), .inData_142(wire_switch_out_stage2[142]), .inData_143(wire_switch_out_stage2[143]), .inData_144(wire_switch_out_stage2[144]), .inData_145(wire_switch_out_stage2[145]), .inData_146(wire_switch_out_stage2[146]), .inData_147(wire_switch_out_stage2[147]), .inData_148(wire_switch_out_stage2[148]), .inData_149(wire_switch_out_stage2[149]), .inData_150(wire_switch_out_stage2[150]), .inData_151(wire_switch_out_stage2[151]), .inData_152(wire_switch_out_stage2[152]), .inData_153(wire_switch_out_stage2[153]), .inData_154(wire_switch_out_stage2[154]), .inData_155(wire_switch_out_stage2[155]), .inData_156(wire_switch_out_stage2[156]), .inData_157(wire_switch_out_stage2[157]), .inData_158(wire_switch_out_stage2[158]), .inData_159(wire_switch_out_stage2[159]), .inData_160(wire_switch_out_stage2[160]), .inData_161(wire_switch_out_stage2[161]), .inData_162(wire_switch_out_stage2[162]), .inData_163(wire_switch_out_stage2[163]), .inData_164(wire_switch_out_stage2[164]), .inData_165(wire_switch_out_stage2[165]), .inData_166(wire_switch_out_stage2[166]), .inData_167(wire_switch_out_stage2[167]), .inData_168(wire_switch_out_stage2[168]), .inData_169(wire_switch_out_stage2[169]), .inData_170(wire_switch_out_stage2[170]), .inData_171(wire_switch_out_stage2[171]), .inData_172(wire_switch_out_stage2[172]), .inData_173(wire_switch_out_stage2[173]), .inData_174(wire_switch_out_stage2[174]), .inData_175(wire_switch_out_stage2[175]), .inData_176(wire_switch_out_stage2[176]), .inData_177(wire_switch_out_stage2[177]), .inData_178(wire_switch_out_stage2[178]), .inData_179(wire_switch_out_stage2[179]), .inData_180(wire_switch_out_stage2[180]), .inData_181(wire_switch_out_stage2[181]), .inData_182(wire_switch_out_stage2[182]), .inData_183(wire_switch_out_stage2[183]), .inData_184(wire_switch_out_stage2[184]), .inData_185(wire_switch_out_stage2[185]), .inData_186(wire_switch_out_stage2[186]), .inData_187(wire_switch_out_stage2[187]), .inData_188(wire_switch_out_stage2[188]), .inData_189(wire_switch_out_stage2[189]), .inData_190(wire_switch_out_stage2[190]), .inData_191(wire_switch_out_stage2[191]), .inData_192(wire_switch_out_stage2[192]), .inData_193(wire_switch_out_stage2[193]), .inData_194(wire_switch_out_stage2[194]), .inData_195(wire_switch_out_stage2[195]), .inData_196(wire_switch_out_stage2[196]), .inData_197(wire_switch_out_stage2[197]), .inData_198(wire_switch_out_stage2[198]), .inData_199(wire_switch_out_stage2[199]), .inData_200(wire_switch_out_stage2[200]), .inData_201(wire_switch_out_stage2[201]), .inData_202(wire_switch_out_stage2[202]), .inData_203(wire_switch_out_stage2[203]), .inData_204(wire_switch_out_stage2[204]), .inData_205(wire_switch_out_stage2[205]), .inData_206(wire_switch_out_stage2[206]), .inData_207(wire_switch_out_stage2[207]), .inData_208(wire_switch_out_stage2[208]), .inData_209(wire_switch_out_stage2[209]), .inData_210(wire_switch_out_stage2[210]), .inData_211(wire_switch_out_stage2[211]), .inData_212(wire_switch_out_stage2[212]), .inData_213(wire_switch_out_stage2[213]), .inData_214(wire_switch_out_stage2[214]), .inData_215(wire_switch_out_stage2[215]), .inData_216(wire_switch_out_stage2[216]), .inData_217(wire_switch_out_stage2[217]), .inData_218(wire_switch_out_stage2[218]), .inData_219(wire_switch_out_stage2[219]), .inData_220(wire_switch_out_stage2[220]), .inData_221(wire_switch_out_stage2[221]), .inData_222(wire_switch_out_stage2[222]), .inData_223(wire_switch_out_stage2[223]), .inData_224(wire_switch_out_stage2[224]), .inData_225(wire_switch_out_stage2[225]), .inData_226(wire_switch_out_stage2[226]), .inData_227(wire_switch_out_stage2[227]), .inData_228(wire_switch_out_stage2[228]), .inData_229(wire_switch_out_stage2[229]), .inData_230(wire_switch_out_stage2[230]), .inData_231(wire_switch_out_stage2[231]), .inData_232(wire_switch_out_stage2[232]), .inData_233(wire_switch_out_stage2[233]), .inData_234(wire_switch_out_stage2[234]), .inData_235(wire_switch_out_stage2[235]), .inData_236(wire_switch_out_stage2[236]), .inData_237(wire_switch_out_stage2[237]), .inData_238(wire_switch_out_stage2[238]), .inData_239(wire_switch_out_stage2[239]), .inData_240(wire_switch_out_stage2[240]), .inData_241(wire_switch_out_stage2[241]), .inData_242(wire_switch_out_stage2[242]), .inData_243(wire_switch_out_stage2[243]), .inData_244(wire_switch_out_stage2[244]), .inData_245(wire_switch_out_stage2[245]), .inData_246(wire_switch_out_stage2[246]), .inData_247(wire_switch_out_stage2[247]), .inData_248(wire_switch_out_stage2[248]), .inData_249(wire_switch_out_stage2[249]), .inData_250(wire_switch_out_stage2[250]), .inData_251(wire_switch_out_stage2[251]), .inData_252(wire_switch_out_stage2[252]), .inData_253(wire_switch_out_stage2[253]), .inData_254(wire_switch_out_stage2[254]), .inData_255(wire_switch_out_stage2[255]), 
        .outData_0(wire_switch_in_stage1[0]), .outData_1(wire_switch_in_stage1[1]), .outData_2(wire_switch_in_stage1[2]), .outData_3(wire_switch_in_stage1[3]), .outData_4(wire_switch_in_stage1[4]), .outData_5(wire_switch_in_stage1[5]), .outData_6(wire_switch_in_stage1[6]), .outData_7(wire_switch_in_stage1[7]), .outData_8(wire_switch_in_stage1[8]), .outData_9(wire_switch_in_stage1[9]), .outData_10(wire_switch_in_stage1[10]), .outData_11(wire_switch_in_stage1[11]), .outData_12(wire_switch_in_stage1[12]), .outData_13(wire_switch_in_stage1[13]), .outData_14(wire_switch_in_stage1[14]), .outData_15(wire_switch_in_stage1[15]), .outData_16(wire_switch_in_stage1[16]), .outData_17(wire_switch_in_stage1[17]), .outData_18(wire_switch_in_stage1[18]), .outData_19(wire_switch_in_stage1[19]), .outData_20(wire_switch_in_stage1[20]), .outData_21(wire_switch_in_stage1[21]), .outData_22(wire_switch_in_stage1[22]), .outData_23(wire_switch_in_stage1[23]), .outData_24(wire_switch_in_stage1[24]), .outData_25(wire_switch_in_stage1[25]), .outData_26(wire_switch_in_stage1[26]), .outData_27(wire_switch_in_stage1[27]), .outData_28(wire_switch_in_stage1[28]), .outData_29(wire_switch_in_stage1[29]), .outData_30(wire_switch_in_stage1[30]), .outData_31(wire_switch_in_stage1[31]), .outData_32(wire_switch_in_stage1[32]), .outData_33(wire_switch_in_stage1[33]), .outData_34(wire_switch_in_stage1[34]), .outData_35(wire_switch_in_stage1[35]), .outData_36(wire_switch_in_stage1[36]), .outData_37(wire_switch_in_stage1[37]), .outData_38(wire_switch_in_stage1[38]), .outData_39(wire_switch_in_stage1[39]), .outData_40(wire_switch_in_stage1[40]), .outData_41(wire_switch_in_stage1[41]), .outData_42(wire_switch_in_stage1[42]), .outData_43(wire_switch_in_stage1[43]), .outData_44(wire_switch_in_stage1[44]), .outData_45(wire_switch_in_stage1[45]), .outData_46(wire_switch_in_stage1[46]), .outData_47(wire_switch_in_stage1[47]), .outData_48(wire_switch_in_stage1[48]), .outData_49(wire_switch_in_stage1[49]), .outData_50(wire_switch_in_stage1[50]), .outData_51(wire_switch_in_stage1[51]), .outData_52(wire_switch_in_stage1[52]), .outData_53(wire_switch_in_stage1[53]), .outData_54(wire_switch_in_stage1[54]), .outData_55(wire_switch_in_stage1[55]), .outData_56(wire_switch_in_stage1[56]), .outData_57(wire_switch_in_stage1[57]), .outData_58(wire_switch_in_stage1[58]), .outData_59(wire_switch_in_stage1[59]), .outData_60(wire_switch_in_stage1[60]), .outData_61(wire_switch_in_stage1[61]), .outData_62(wire_switch_in_stage1[62]), .outData_63(wire_switch_in_stage1[63]), .outData_64(wire_switch_in_stage1[64]), .outData_65(wire_switch_in_stage1[65]), .outData_66(wire_switch_in_stage1[66]), .outData_67(wire_switch_in_stage1[67]), .outData_68(wire_switch_in_stage1[68]), .outData_69(wire_switch_in_stage1[69]), .outData_70(wire_switch_in_stage1[70]), .outData_71(wire_switch_in_stage1[71]), .outData_72(wire_switch_in_stage1[72]), .outData_73(wire_switch_in_stage1[73]), .outData_74(wire_switch_in_stage1[74]), .outData_75(wire_switch_in_stage1[75]), .outData_76(wire_switch_in_stage1[76]), .outData_77(wire_switch_in_stage1[77]), .outData_78(wire_switch_in_stage1[78]), .outData_79(wire_switch_in_stage1[79]), .outData_80(wire_switch_in_stage1[80]), .outData_81(wire_switch_in_stage1[81]), .outData_82(wire_switch_in_stage1[82]), .outData_83(wire_switch_in_stage1[83]), .outData_84(wire_switch_in_stage1[84]), .outData_85(wire_switch_in_stage1[85]), .outData_86(wire_switch_in_stage1[86]), .outData_87(wire_switch_in_stage1[87]), .outData_88(wire_switch_in_stage1[88]), .outData_89(wire_switch_in_stage1[89]), .outData_90(wire_switch_in_stage1[90]), .outData_91(wire_switch_in_stage1[91]), .outData_92(wire_switch_in_stage1[92]), .outData_93(wire_switch_in_stage1[93]), .outData_94(wire_switch_in_stage1[94]), .outData_95(wire_switch_in_stage1[95]), .outData_96(wire_switch_in_stage1[96]), .outData_97(wire_switch_in_stage1[97]), .outData_98(wire_switch_in_stage1[98]), .outData_99(wire_switch_in_stage1[99]), .outData_100(wire_switch_in_stage1[100]), .outData_101(wire_switch_in_stage1[101]), .outData_102(wire_switch_in_stage1[102]), .outData_103(wire_switch_in_stage1[103]), .outData_104(wire_switch_in_stage1[104]), .outData_105(wire_switch_in_stage1[105]), .outData_106(wire_switch_in_stage1[106]), .outData_107(wire_switch_in_stage1[107]), .outData_108(wire_switch_in_stage1[108]), .outData_109(wire_switch_in_stage1[109]), .outData_110(wire_switch_in_stage1[110]), .outData_111(wire_switch_in_stage1[111]), .outData_112(wire_switch_in_stage1[112]), .outData_113(wire_switch_in_stage1[113]), .outData_114(wire_switch_in_stage1[114]), .outData_115(wire_switch_in_stage1[115]), .outData_116(wire_switch_in_stage1[116]), .outData_117(wire_switch_in_stage1[117]), .outData_118(wire_switch_in_stage1[118]), .outData_119(wire_switch_in_stage1[119]), .outData_120(wire_switch_in_stage1[120]), .outData_121(wire_switch_in_stage1[121]), .outData_122(wire_switch_in_stage1[122]), .outData_123(wire_switch_in_stage1[123]), .outData_124(wire_switch_in_stage1[124]), .outData_125(wire_switch_in_stage1[125]), .outData_126(wire_switch_in_stage1[126]), .outData_127(wire_switch_in_stage1[127]), .outData_128(wire_switch_in_stage1[128]), .outData_129(wire_switch_in_stage1[129]), .outData_130(wire_switch_in_stage1[130]), .outData_131(wire_switch_in_stage1[131]), .outData_132(wire_switch_in_stage1[132]), .outData_133(wire_switch_in_stage1[133]), .outData_134(wire_switch_in_stage1[134]), .outData_135(wire_switch_in_stage1[135]), .outData_136(wire_switch_in_stage1[136]), .outData_137(wire_switch_in_stage1[137]), .outData_138(wire_switch_in_stage1[138]), .outData_139(wire_switch_in_stage1[139]), .outData_140(wire_switch_in_stage1[140]), .outData_141(wire_switch_in_stage1[141]), .outData_142(wire_switch_in_stage1[142]), .outData_143(wire_switch_in_stage1[143]), .outData_144(wire_switch_in_stage1[144]), .outData_145(wire_switch_in_stage1[145]), .outData_146(wire_switch_in_stage1[146]), .outData_147(wire_switch_in_stage1[147]), .outData_148(wire_switch_in_stage1[148]), .outData_149(wire_switch_in_stage1[149]), .outData_150(wire_switch_in_stage1[150]), .outData_151(wire_switch_in_stage1[151]), .outData_152(wire_switch_in_stage1[152]), .outData_153(wire_switch_in_stage1[153]), .outData_154(wire_switch_in_stage1[154]), .outData_155(wire_switch_in_stage1[155]), .outData_156(wire_switch_in_stage1[156]), .outData_157(wire_switch_in_stage1[157]), .outData_158(wire_switch_in_stage1[158]), .outData_159(wire_switch_in_stage1[159]), .outData_160(wire_switch_in_stage1[160]), .outData_161(wire_switch_in_stage1[161]), .outData_162(wire_switch_in_stage1[162]), .outData_163(wire_switch_in_stage1[163]), .outData_164(wire_switch_in_stage1[164]), .outData_165(wire_switch_in_stage1[165]), .outData_166(wire_switch_in_stage1[166]), .outData_167(wire_switch_in_stage1[167]), .outData_168(wire_switch_in_stage1[168]), .outData_169(wire_switch_in_stage1[169]), .outData_170(wire_switch_in_stage1[170]), .outData_171(wire_switch_in_stage1[171]), .outData_172(wire_switch_in_stage1[172]), .outData_173(wire_switch_in_stage1[173]), .outData_174(wire_switch_in_stage1[174]), .outData_175(wire_switch_in_stage1[175]), .outData_176(wire_switch_in_stage1[176]), .outData_177(wire_switch_in_stage1[177]), .outData_178(wire_switch_in_stage1[178]), .outData_179(wire_switch_in_stage1[179]), .outData_180(wire_switch_in_stage1[180]), .outData_181(wire_switch_in_stage1[181]), .outData_182(wire_switch_in_stage1[182]), .outData_183(wire_switch_in_stage1[183]), .outData_184(wire_switch_in_stage1[184]), .outData_185(wire_switch_in_stage1[185]), .outData_186(wire_switch_in_stage1[186]), .outData_187(wire_switch_in_stage1[187]), .outData_188(wire_switch_in_stage1[188]), .outData_189(wire_switch_in_stage1[189]), .outData_190(wire_switch_in_stage1[190]), .outData_191(wire_switch_in_stage1[191]), .outData_192(wire_switch_in_stage1[192]), .outData_193(wire_switch_in_stage1[193]), .outData_194(wire_switch_in_stage1[194]), .outData_195(wire_switch_in_stage1[195]), .outData_196(wire_switch_in_stage1[196]), .outData_197(wire_switch_in_stage1[197]), .outData_198(wire_switch_in_stage1[198]), .outData_199(wire_switch_in_stage1[199]), .outData_200(wire_switch_in_stage1[200]), .outData_201(wire_switch_in_stage1[201]), .outData_202(wire_switch_in_stage1[202]), .outData_203(wire_switch_in_stage1[203]), .outData_204(wire_switch_in_stage1[204]), .outData_205(wire_switch_in_stage1[205]), .outData_206(wire_switch_in_stage1[206]), .outData_207(wire_switch_in_stage1[207]), .outData_208(wire_switch_in_stage1[208]), .outData_209(wire_switch_in_stage1[209]), .outData_210(wire_switch_in_stage1[210]), .outData_211(wire_switch_in_stage1[211]), .outData_212(wire_switch_in_stage1[212]), .outData_213(wire_switch_in_stage1[213]), .outData_214(wire_switch_in_stage1[214]), .outData_215(wire_switch_in_stage1[215]), .outData_216(wire_switch_in_stage1[216]), .outData_217(wire_switch_in_stage1[217]), .outData_218(wire_switch_in_stage1[218]), .outData_219(wire_switch_in_stage1[219]), .outData_220(wire_switch_in_stage1[220]), .outData_221(wire_switch_in_stage1[221]), .outData_222(wire_switch_in_stage1[222]), .outData_223(wire_switch_in_stage1[223]), .outData_224(wire_switch_in_stage1[224]), .outData_225(wire_switch_in_stage1[225]), .outData_226(wire_switch_in_stage1[226]), .outData_227(wire_switch_in_stage1[227]), .outData_228(wire_switch_in_stage1[228]), .outData_229(wire_switch_in_stage1[229]), .outData_230(wire_switch_in_stage1[230]), .outData_231(wire_switch_in_stage1[231]), .outData_232(wire_switch_in_stage1[232]), .outData_233(wire_switch_in_stage1[233]), .outData_234(wire_switch_in_stage1[234]), .outData_235(wire_switch_in_stage1[235]), .outData_236(wire_switch_in_stage1[236]), .outData_237(wire_switch_in_stage1[237]), .outData_238(wire_switch_in_stage1[238]), .outData_239(wire_switch_in_stage1[239]), .outData_240(wire_switch_in_stage1[240]), .outData_241(wire_switch_in_stage1[241]), .outData_242(wire_switch_in_stage1[242]), .outData_243(wire_switch_in_stage1[243]), .outData_244(wire_switch_in_stage1[244]), .outData_245(wire_switch_in_stage1[245]), .outData_246(wire_switch_in_stage1[246]), .outData_247(wire_switch_in_stage1[247]), .outData_248(wire_switch_in_stage1[248]), .outData_249(wire_switch_in_stage1[249]), .outData_250(wire_switch_in_stage1[250]), .outData_251(wire_switch_in_stage1[251]), .outData_252(wire_switch_in_stage1[252]), .outData_253(wire_switch_in_stage1[253]), .outData_254(wire_switch_in_stage1[254]), .outData_255(wire_switch_in_stage1[255]), 
        .in_start(in_start_stage1), .out_start(con_in_start_stage1), .clk(clk), .rst(rst)); 

  
  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[0] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[1] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[2] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[3] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[4] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[5] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[6] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[7] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[8] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[9] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[10] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[11] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[12] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[13] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[14] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[15] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[16] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[17] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[18] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[19] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[20] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[21] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[22] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[23] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[24] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[25] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[26] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[27] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[28] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[29] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[30] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[31] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[32] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[33] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[34] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[35] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[36] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[37] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[38] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[39] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[40] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[41] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[42] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[43] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[44] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[45] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[46] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[47] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[48] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[49] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[50] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[51] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[52] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[53] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[54] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[55] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[56] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[57] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[58] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[59] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[60] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[61] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[62] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[63] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[64] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[65] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[66] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[67] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[68] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[69] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[70] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[71] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[72] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[73] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[74] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[75] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[76] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[77] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[78] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[79] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[80] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[81] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[82] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[83] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[84] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[85] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[86] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[87] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[88] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[89] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[90] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[91] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[92] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[93] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[94] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[95] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[96] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[97] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[98] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[99] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[100] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[101] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[102] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[103] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[104] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[105] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[106] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[107] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[108] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[109] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[110] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[111] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[112] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[113] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[114] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[115] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[116] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[117] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[118] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[119] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[120] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[121] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[122] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[123] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[124] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[125] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[126] <= counter_w[6]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage1[127] <= counter_w[6]; 
  end                            

  wire [DATA_WIDTH-1:0] wire_switch_in_stage0[255:0];
  wire [DATA_WIDTH-1:0] wire_switch_out_stage0[255:0];
  reg [127:0] wire_ctrl_stage0;

  switches_stage_st0_0_R switch_stage_0(
        .inData_0(wire_switch_in_stage0[0]), .inData_1(wire_switch_in_stage0[1]), .inData_2(wire_switch_in_stage0[2]), .inData_3(wire_switch_in_stage0[3]), .inData_4(wire_switch_in_stage0[4]), .inData_5(wire_switch_in_stage0[5]), .inData_6(wire_switch_in_stage0[6]), .inData_7(wire_switch_in_stage0[7]), .inData_8(wire_switch_in_stage0[8]), .inData_9(wire_switch_in_stage0[9]), .inData_10(wire_switch_in_stage0[10]), .inData_11(wire_switch_in_stage0[11]), .inData_12(wire_switch_in_stage0[12]), .inData_13(wire_switch_in_stage0[13]), .inData_14(wire_switch_in_stage0[14]), .inData_15(wire_switch_in_stage0[15]), .inData_16(wire_switch_in_stage0[16]), .inData_17(wire_switch_in_stage0[17]), .inData_18(wire_switch_in_stage0[18]), .inData_19(wire_switch_in_stage0[19]), .inData_20(wire_switch_in_stage0[20]), .inData_21(wire_switch_in_stage0[21]), .inData_22(wire_switch_in_stage0[22]), .inData_23(wire_switch_in_stage0[23]), .inData_24(wire_switch_in_stage0[24]), .inData_25(wire_switch_in_stage0[25]), .inData_26(wire_switch_in_stage0[26]), .inData_27(wire_switch_in_stage0[27]), .inData_28(wire_switch_in_stage0[28]), .inData_29(wire_switch_in_stage0[29]), .inData_30(wire_switch_in_stage0[30]), .inData_31(wire_switch_in_stage0[31]), .inData_32(wire_switch_in_stage0[32]), .inData_33(wire_switch_in_stage0[33]), .inData_34(wire_switch_in_stage0[34]), .inData_35(wire_switch_in_stage0[35]), .inData_36(wire_switch_in_stage0[36]), .inData_37(wire_switch_in_stage0[37]), .inData_38(wire_switch_in_stage0[38]), .inData_39(wire_switch_in_stage0[39]), .inData_40(wire_switch_in_stage0[40]), .inData_41(wire_switch_in_stage0[41]), .inData_42(wire_switch_in_stage0[42]), .inData_43(wire_switch_in_stage0[43]), .inData_44(wire_switch_in_stage0[44]), .inData_45(wire_switch_in_stage0[45]), .inData_46(wire_switch_in_stage0[46]), .inData_47(wire_switch_in_stage0[47]), .inData_48(wire_switch_in_stage0[48]), .inData_49(wire_switch_in_stage0[49]), .inData_50(wire_switch_in_stage0[50]), .inData_51(wire_switch_in_stage0[51]), .inData_52(wire_switch_in_stage0[52]), .inData_53(wire_switch_in_stage0[53]), .inData_54(wire_switch_in_stage0[54]), .inData_55(wire_switch_in_stage0[55]), .inData_56(wire_switch_in_stage0[56]), .inData_57(wire_switch_in_stage0[57]), .inData_58(wire_switch_in_stage0[58]), .inData_59(wire_switch_in_stage0[59]), .inData_60(wire_switch_in_stage0[60]), .inData_61(wire_switch_in_stage0[61]), .inData_62(wire_switch_in_stage0[62]), .inData_63(wire_switch_in_stage0[63]), .inData_64(wire_switch_in_stage0[64]), .inData_65(wire_switch_in_stage0[65]), .inData_66(wire_switch_in_stage0[66]), .inData_67(wire_switch_in_stage0[67]), .inData_68(wire_switch_in_stage0[68]), .inData_69(wire_switch_in_stage0[69]), .inData_70(wire_switch_in_stage0[70]), .inData_71(wire_switch_in_stage0[71]), .inData_72(wire_switch_in_stage0[72]), .inData_73(wire_switch_in_stage0[73]), .inData_74(wire_switch_in_stage0[74]), .inData_75(wire_switch_in_stage0[75]), .inData_76(wire_switch_in_stage0[76]), .inData_77(wire_switch_in_stage0[77]), .inData_78(wire_switch_in_stage0[78]), .inData_79(wire_switch_in_stage0[79]), .inData_80(wire_switch_in_stage0[80]), .inData_81(wire_switch_in_stage0[81]), .inData_82(wire_switch_in_stage0[82]), .inData_83(wire_switch_in_stage0[83]), .inData_84(wire_switch_in_stage0[84]), .inData_85(wire_switch_in_stage0[85]), .inData_86(wire_switch_in_stage0[86]), .inData_87(wire_switch_in_stage0[87]), .inData_88(wire_switch_in_stage0[88]), .inData_89(wire_switch_in_stage0[89]), .inData_90(wire_switch_in_stage0[90]), .inData_91(wire_switch_in_stage0[91]), .inData_92(wire_switch_in_stage0[92]), .inData_93(wire_switch_in_stage0[93]), .inData_94(wire_switch_in_stage0[94]), .inData_95(wire_switch_in_stage0[95]), .inData_96(wire_switch_in_stage0[96]), .inData_97(wire_switch_in_stage0[97]), .inData_98(wire_switch_in_stage0[98]), .inData_99(wire_switch_in_stage0[99]), .inData_100(wire_switch_in_stage0[100]), .inData_101(wire_switch_in_stage0[101]), .inData_102(wire_switch_in_stage0[102]), .inData_103(wire_switch_in_stage0[103]), .inData_104(wire_switch_in_stage0[104]), .inData_105(wire_switch_in_stage0[105]), .inData_106(wire_switch_in_stage0[106]), .inData_107(wire_switch_in_stage0[107]), .inData_108(wire_switch_in_stage0[108]), .inData_109(wire_switch_in_stage0[109]), .inData_110(wire_switch_in_stage0[110]), .inData_111(wire_switch_in_stage0[111]), .inData_112(wire_switch_in_stage0[112]), .inData_113(wire_switch_in_stage0[113]), .inData_114(wire_switch_in_stage0[114]), .inData_115(wire_switch_in_stage0[115]), .inData_116(wire_switch_in_stage0[116]), .inData_117(wire_switch_in_stage0[117]), .inData_118(wire_switch_in_stage0[118]), .inData_119(wire_switch_in_stage0[119]), .inData_120(wire_switch_in_stage0[120]), .inData_121(wire_switch_in_stage0[121]), .inData_122(wire_switch_in_stage0[122]), .inData_123(wire_switch_in_stage0[123]), .inData_124(wire_switch_in_stage0[124]), .inData_125(wire_switch_in_stage0[125]), .inData_126(wire_switch_in_stage0[126]), .inData_127(wire_switch_in_stage0[127]), .inData_128(wire_switch_in_stage0[128]), .inData_129(wire_switch_in_stage0[129]), .inData_130(wire_switch_in_stage0[130]), .inData_131(wire_switch_in_stage0[131]), .inData_132(wire_switch_in_stage0[132]), .inData_133(wire_switch_in_stage0[133]), .inData_134(wire_switch_in_stage0[134]), .inData_135(wire_switch_in_stage0[135]), .inData_136(wire_switch_in_stage0[136]), .inData_137(wire_switch_in_stage0[137]), .inData_138(wire_switch_in_stage0[138]), .inData_139(wire_switch_in_stage0[139]), .inData_140(wire_switch_in_stage0[140]), .inData_141(wire_switch_in_stage0[141]), .inData_142(wire_switch_in_stage0[142]), .inData_143(wire_switch_in_stage0[143]), .inData_144(wire_switch_in_stage0[144]), .inData_145(wire_switch_in_stage0[145]), .inData_146(wire_switch_in_stage0[146]), .inData_147(wire_switch_in_stage0[147]), .inData_148(wire_switch_in_stage0[148]), .inData_149(wire_switch_in_stage0[149]), .inData_150(wire_switch_in_stage0[150]), .inData_151(wire_switch_in_stage0[151]), .inData_152(wire_switch_in_stage0[152]), .inData_153(wire_switch_in_stage0[153]), .inData_154(wire_switch_in_stage0[154]), .inData_155(wire_switch_in_stage0[155]), .inData_156(wire_switch_in_stage0[156]), .inData_157(wire_switch_in_stage0[157]), .inData_158(wire_switch_in_stage0[158]), .inData_159(wire_switch_in_stage0[159]), .inData_160(wire_switch_in_stage0[160]), .inData_161(wire_switch_in_stage0[161]), .inData_162(wire_switch_in_stage0[162]), .inData_163(wire_switch_in_stage0[163]), .inData_164(wire_switch_in_stage0[164]), .inData_165(wire_switch_in_stage0[165]), .inData_166(wire_switch_in_stage0[166]), .inData_167(wire_switch_in_stage0[167]), .inData_168(wire_switch_in_stage0[168]), .inData_169(wire_switch_in_stage0[169]), .inData_170(wire_switch_in_stage0[170]), .inData_171(wire_switch_in_stage0[171]), .inData_172(wire_switch_in_stage0[172]), .inData_173(wire_switch_in_stage0[173]), .inData_174(wire_switch_in_stage0[174]), .inData_175(wire_switch_in_stage0[175]), .inData_176(wire_switch_in_stage0[176]), .inData_177(wire_switch_in_stage0[177]), .inData_178(wire_switch_in_stage0[178]), .inData_179(wire_switch_in_stage0[179]), .inData_180(wire_switch_in_stage0[180]), .inData_181(wire_switch_in_stage0[181]), .inData_182(wire_switch_in_stage0[182]), .inData_183(wire_switch_in_stage0[183]), .inData_184(wire_switch_in_stage0[184]), .inData_185(wire_switch_in_stage0[185]), .inData_186(wire_switch_in_stage0[186]), .inData_187(wire_switch_in_stage0[187]), .inData_188(wire_switch_in_stage0[188]), .inData_189(wire_switch_in_stage0[189]), .inData_190(wire_switch_in_stage0[190]), .inData_191(wire_switch_in_stage0[191]), .inData_192(wire_switch_in_stage0[192]), .inData_193(wire_switch_in_stage0[193]), .inData_194(wire_switch_in_stage0[194]), .inData_195(wire_switch_in_stage0[195]), .inData_196(wire_switch_in_stage0[196]), .inData_197(wire_switch_in_stage0[197]), .inData_198(wire_switch_in_stage0[198]), .inData_199(wire_switch_in_stage0[199]), .inData_200(wire_switch_in_stage0[200]), .inData_201(wire_switch_in_stage0[201]), .inData_202(wire_switch_in_stage0[202]), .inData_203(wire_switch_in_stage0[203]), .inData_204(wire_switch_in_stage0[204]), .inData_205(wire_switch_in_stage0[205]), .inData_206(wire_switch_in_stage0[206]), .inData_207(wire_switch_in_stage0[207]), .inData_208(wire_switch_in_stage0[208]), .inData_209(wire_switch_in_stage0[209]), .inData_210(wire_switch_in_stage0[210]), .inData_211(wire_switch_in_stage0[211]), .inData_212(wire_switch_in_stage0[212]), .inData_213(wire_switch_in_stage0[213]), .inData_214(wire_switch_in_stage0[214]), .inData_215(wire_switch_in_stage0[215]), .inData_216(wire_switch_in_stage0[216]), .inData_217(wire_switch_in_stage0[217]), .inData_218(wire_switch_in_stage0[218]), .inData_219(wire_switch_in_stage0[219]), .inData_220(wire_switch_in_stage0[220]), .inData_221(wire_switch_in_stage0[221]), .inData_222(wire_switch_in_stage0[222]), .inData_223(wire_switch_in_stage0[223]), .inData_224(wire_switch_in_stage0[224]), .inData_225(wire_switch_in_stage0[225]), .inData_226(wire_switch_in_stage0[226]), .inData_227(wire_switch_in_stage0[227]), .inData_228(wire_switch_in_stage0[228]), .inData_229(wire_switch_in_stage0[229]), .inData_230(wire_switch_in_stage0[230]), .inData_231(wire_switch_in_stage0[231]), .inData_232(wire_switch_in_stage0[232]), .inData_233(wire_switch_in_stage0[233]), .inData_234(wire_switch_in_stage0[234]), .inData_235(wire_switch_in_stage0[235]), .inData_236(wire_switch_in_stage0[236]), .inData_237(wire_switch_in_stage0[237]), .inData_238(wire_switch_in_stage0[238]), .inData_239(wire_switch_in_stage0[239]), .inData_240(wire_switch_in_stage0[240]), .inData_241(wire_switch_in_stage0[241]), .inData_242(wire_switch_in_stage0[242]), .inData_243(wire_switch_in_stage0[243]), .inData_244(wire_switch_in_stage0[244]), .inData_245(wire_switch_in_stage0[245]), .inData_246(wire_switch_in_stage0[246]), .inData_247(wire_switch_in_stage0[247]), .inData_248(wire_switch_in_stage0[248]), .inData_249(wire_switch_in_stage0[249]), .inData_250(wire_switch_in_stage0[250]), .inData_251(wire_switch_in_stage0[251]), .inData_252(wire_switch_in_stage0[252]), .inData_253(wire_switch_in_stage0[253]), .inData_254(wire_switch_in_stage0[254]), .inData_255(wire_switch_in_stage0[255]), 
        .outData_0(wireOut[0]), .outData_1(wireOut[1]), .outData_2(wireOut[2]), .outData_3(wireOut[3]), .outData_4(wireOut[4]), .outData_5(wireOut[5]), .outData_6(wireOut[6]), .outData_7(wireOut[7]), .outData_8(wireOut[8]), .outData_9(wireOut[9]), .outData_10(wireOut[10]), .outData_11(wireOut[11]), .outData_12(wireOut[12]), .outData_13(wireOut[13]), .outData_14(wireOut[14]), .outData_15(wireOut[15]), .outData_16(wireOut[16]), .outData_17(wireOut[17]), .outData_18(wireOut[18]), .outData_19(wireOut[19]), .outData_20(wireOut[20]), .outData_21(wireOut[21]), .outData_22(wireOut[22]), .outData_23(wireOut[23]), .outData_24(wireOut[24]), .outData_25(wireOut[25]), .outData_26(wireOut[26]), .outData_27(wireOut[27]), .outData_28(wireOut[28]), .outData_29(wireOut[29]), .outData_30(wireOut[30]), .outData_31(wireOut[31]), .outData_32(wireOut[32]), .outData_33(wireOut[33]), .outData_34(wireOut[34]), .outData_35(wireOut[35]), .outData_36(wireOut[36]), .outData_37(wireOut[37]), .outData_38(wireOut[38]), .outData_39(wireOut[39]), .outData_40(wireOut[40]), .outData_41(wireOut[41]), .outData_42(wireOut[42]), .outData_43(wireOut[43]), .outData_44(wireOut[44]), .outData_45(wireOut[45]), .outData_46(wireOut[46]), .outData_47(wireOut[47]), .outData_48(wireOut[48]), .outData_49(wireOut[49]), .outData_50(wireOut[50]), .outData_51(wireOut[51]), .outData_52(wireOut[52]), .outData_53(wireOut[53]), .outData_54(wireOut[54]), .outData_55(wireOut[55]), .outData_56(wireOut[56]), .outData_57(wireOut[57]), .outData_58(wireOut[58]), .outData_59(wireOut[59]), .outData_60(wireOut[60]), .outData_61(wireOut[61]), .outData_62(wireOut[62]), .outData_63(wireOut[63]), .outData_64(wireOut[64]), .outData_65(wireOut[65]), .outData_66(wireOut[66]), .outData_67(wireOut[67]), .outData_68(wireOut[68]), .outData_69(wireOut[69]), .outData_70(wireOut[70]), .outData_71(wireOut[71]), .outData_72(wireOut[72]), .outData_73(wireOut[73]), .outData_74(wireOut[74]), .outData_75(wireOut[75]), .outData_76(wireOut[76]), .outData_77(wireOut[77]), .outData_78(wireOut[78]), .outData_79(wireOut[79]), .outData_80(wireOut[80]), .outData_81(wireOut[81]), .outData_82(wireOut[82]), .outData_83(wireOut[83]), .outData_84(wireOut[84]), .outData_85(wireOut[85]), .outData_86(wireOut[86]), .outData_87(wireOut[87]), .outData_88(wireOut[88]), .outData_89(wireOut[89]), .outData_90(wireOut[90]), .outData_91(wireOut[91]), .outData_92(wireOut[92]), .outData_93(wireOut[93]), .outData_94(wireOut[94]), .outData_95(wireOut[95]), .outData_96(wireOut[96]), .outData_97(wireOut[97]), .outData_98(wireOut[98]), .outData_99(wireOut[99]), .outData_100(wireOut[100]), .outData_101(wireOut[101]), .outData_102(wireOut[102]), .outData_103(wireOut[103]), .outData_104(wireOut[104]), .outData_105(wireOut[105]), .outData_106(wireOut[106]), .outData_107(wireOut[107]), .outData_108(wireOut[108]), .outData_109(wireOut[109]), .outData_110(wireOut[110]), .outData_111(wireOut[111]), .outData_112(wireOut[112]), .outData_113(wireOut[113]), .outData_114(wireOut[114]), .outData_115(wireOut[115]), .outData_116(wireOut[116]), .outData_117(wireOut[117]), .outData_118(wireOut[118]), .outData_119(wireOut[119]), .outData_120(wireOut[120]), .outData_121(wireOut[121]), .outData_122(wireOut[122]), .outData_123(wireOut[123]), .outData_124(wireOut[124]), .outData_125(wireOut[125]), .outData_126(wireOut[126]), .outData_127(wireOut[127]), .outData_128(wireOut[128]), .outData_129(wireOut[129]), .outData_130(wireOut[130]), .outData_131(wireOut[131]), .outData_132(wireOut[132]), .outData_133(wireOut[133]), .outData_134(wireOut[134]), .outData_135(wireOut[135]), .outData_136(wireOut[136]), .outData_137(wireOut[137]), .outData_138(wireOut[138]), .outData_139(wireOut[139]), .outData_140(wireOut[140]), .outData_141(wireOut[141]), .outData_142(wireOut[142]), .outData_143(wireOut[143]), .outData_144(wireOut[144]), .outData_145(wireOut[145]), .outData_146(wireOut[146]), .outData_147(wireOut[147]), .outData_148(wireOut[148]), .outData_149(wireOut[149]), .outData_150(wireOut[150]), .outData_151(wireOut[151]), .outData_152(wireOut[152]), .outData_153(wireOut[153]), .outData_154(wireOut[154]), .outData_155(wireOut[155]), .outData_156(wireOut[156]), .outData_157(wireOut[157]), .outData_158(wireOut[158]), .outData_159(wireOut[159]), .outData_160(wireOut[160]), .outData_161(wireOut[161]), .outData_162(wireOut[162]), .outData_163(wireOut[163]), .outData_164(wireOut[164]), .outData_165(wireOut[165]), .outData_166(wireOut[166]), .outData_167(wireOut[167]), .outData_168(wireOut[168]), .outData_169(wireOut[169]), .outData_170(wireOut[170]), .outData_171(wireOut[171]), .outData_172(wireOut[172]), .outData_173(wireOut[173]), .outData_174(wireOut[174]), .outData_175(wireOut[175]), .outData_176(wireOut[176]), .outData_177(wireOut[177]), .outData_178(wireOut[178]), .outData_179(wireOut[179]), .outData_180(wireOut[180]), .outData_181(wireOut[181]), .outData_182(wireOut[182]), .outData_183(wireOut[183]), .outData_184(wireOut[184]), .outData_185(wireOut[185]), .outData_186(wireOut[186]), .outData_187(wireOut[187]), .outData_188(wireOut[188]), .outData_189(wireOut[189]), .outData_190(wireOut[190]), .outData_191(wireOut[191]), .outData_192(wireOut[192]), .outData_193(wireOut[193]), .outData_194(wireOut[194]), .outData_195(wireOut[195]), .outData_196(wireOut[196]), .outData_197(wireOut[197]), .outData_198(wireOut[198]), .outData_199(wireOut[199]), .outData_200(wireOut[200]), .outData_201(wireOut[201]), .outData_202(wireOut[202]), .outData_203(wireOut[203]), .outData_204(wireOut[204]), .outData_205(wireOut[205]), .outData_206(wireOut[206]), .outData_207(wireOut[207]), .outData_208(wireOut[208]), .outData_209(wireOut[209]), .outData_210(wireOut[210]), .outData_211(wireOut[211]), .outData_212(wireOut[212]), .outData_213(wireOut[213]), .outData_214(wireOut[214]), .outData_215(wireOut[215]), .outData_216(wireOut[216]), .outData_217(wireOut[217]), .outData_218(wireOut[218]), .outData_219(wireOut[219]), .outData_220(wireOut[220]), .outData_221(wireOut[221]), .outData_222(wireOut[222]), .outData_223(wireOut[223]), .outData_224(wireOut[224]), .outData_225(wireOut[225]), .outData_226(wireOut[226]), .outData_227(wireOut[227]), .outData_228(wireOut[228]), .outData_229(wireOut[229]), .outData_230(wireOut[230]), .outData_231(wireOut[231]), .outData_232(wireOut[232]), .outData_233(wireOut[233]), .outData_234(wireOut[234]), .outData_235(wireOut[235]), .outData_236(wireOut[236]), .outData_237(wireOut[237]), .outData_238(wireOut[238]), .outData_239(wireOut[239]), .outData_240(wireOut[240]), .outData_241(wireOut[241]), .outData_242(wireOut[242]), .outData_243(wireOut[243]), .outData_244(wireOut[244]), .outData_245(wireOut[245]), .outData_246(wireOut[246]), .outData_247(wireOut[247]), .outData_248(wireOut[248]), .outData_249(wireOut[249]), .outData_250(wireOut[250]), .outData_251(wireOut[251]), .outData_252(wireOut[252]), .outData_253(wireOut[253]), .outData_254(wireOut[254]), .outData_255(wireOut[255]), 
        .in_start(con_in_start_stage0), .out_start(out_start_w), .ctrl(wire_ctrl_stage0), .clk(clk), .rst(rst));
  
  wireCon_dp256_st0_R wire_stage_0(
        .inData_0(wire_switch_out_stage1[0]), .inData_1(wire_switch_out_stage1[1]), .inData_2(wire_switch_out_stage1[2]), .inData_3(wire_switch_out_stage1[3]), .inData_4(wire_switch_out_stage1[4]), .inData_5(wire_switch_out_stage1[5]), .inData_6(wire_switch_out_stage1[6]), .inData_7(wire_switch_out_stage1[7]), .inData_8(wire_switch_out_stage1[8]), .inData_9(wire_switch_out_stage1[9]), .inData_10(wire_switch_out_stage1[10]), .inData_11(wire_switch_out_stage1[11]), .inData_12(wire_switch_out_stage1[12]), .inData_13(wire_switch_out_stage1[13]), .inData_14(wire_switch_out_stage1[14]), .inData_15(wire_switch_out_stage1[15]), .inData_16(wire_switch_out_stage1[16]), .inData_17(wire_switch_out_stage1[17]), .inData_18(wire_switch_out_stage1[18]), .inData_19(wire_switch_out_stage1[19]), .inData_20(wire_switch_out_stage1[20]), .inData_21(wire_switch_out_stage1[21]), .inData_22(wire_switch_out_stage1[22]), .inData_23(wire_switch_out_stage1[23]), .inData_24(wire_switch_out_stage1[24]), .inData_25(wire_switch_out_stage1[25]), .inData_26(wire_switch_out_stage1[26]), .inData_27(wire_switch_out_stage1[27]), .inData_28(wire_switch_out_stage1[28]), .inData_29(wire_switch_out_stage1[29]), .inData_30(wire_switch_out_stage1[30]), .inData_31(wire_switch_out_stage1[31]), .inData_32(wire_switch_out_stage1[32]), .inData_33(wire_switch_out_stage1[33]), .inData_34(wire_switch_out_stage1[34]), .inData_35(wire_switch_out_stage1[35]), .inData_36(wire_switch_out_stage1[36]), .inData_37(wire_switch_out_stage1[37]), .inData_38(wire_switch_out_stage1[38]), .inData_39(wire_switch_out_stage1[39]), .inData_40(wire_switch_out_stage1[40]), .inData_41(wire_switch_out_stage1[41]), .inData_42(wire_switch_out_stage1[42]), .inData_43(wire_switch_out_stage1[43]), .inData_44(wire_switch_out_stage1[44]), .inData_45(wire_switch_out_stage1[45]), .inData_46(wire_switch_out_stage1[46]), .inData_47(wire_switch_out_stage1[47]), .inData_48(wire_switch_out_stage1[48]), .inData_49(wire_switch_out_stage1[49]), .inData_50(wire_switch_out_stage1[50]), .inData_51(wire_switch_out_stage1[51]), .inData_52(wire_switch_out_stage1[52]), .inData_53(wire_switch_out_stage1[53]), .inData_54(wire_switch_out_stage1[54]), .inData_55(wire_switch_out_stage1[55]), .inData_56(wire_switch_out_stage1[56]), .inData_57(wire_switch_out_stage1[57]), .inData_58(wire_switch_out_stage1[58]), .inData_59(wire_switch_out_stage1[59]), .inData_60(wire_switch_out_stage1[60]), .inData_61(wire_switch_out_stage1[61]), .inData_62(wire_switch_out_stage1[62]), .inData_63(wire_switch_out_stage1[63]), .inData_64(wire_switch_out_stage1[64]), .inData_65(wire_switch_out_stage1[65]), .inData_66(wire_switch_out_stage1[66]), .inData_67(wire_switch_out_stage1[67]), .inData_68(wire_switch_out_stage1[68]), .inData_69(wire_switch_out_stage1[69]), .inData_70(wire_switch_out_stage1[70]), .inData_71(wire_switch_out_stage1[71]), .inData_72(wire_switch_out_stage1[72]), .inData_73(wire_switch_out_stage1[73]), .inData_74(wire_switch_out_stage1[74]), .inData_75(wire_switch_out_stage1[75]), .inData_76(wire_switch_out_stage1[76]), .inData_77(wire_switch_out_stage1[77]), .inData_78(wire_switch_out_stage1[78]), .inData_79(wire_switch_out_stage1[79]), .inData_80(wire_switch_out_stage1[80]), .inData_81(wire_switch_out_stage1[81]), .inData_82(wire_switch_out_stage1[82]), .inData_83(wire_switch_out_stage1[83]), .inData_84(wire_switch_out_stage1[84]), .inData_85(wire_switch_out_stage1[85]), .inData_86(wire_switch_out_stage1[86]), .inData_87(wire_switch_out_stage1[87]), .inData_88(wire_switch_out_stage1[88]), .inData_89(wire_switch_out_stage1[89]), .inData_90(wire_switch_out_stage1[90]), .inData_91(wire_switch_out_stage1[91]), .inData_92(wire_switch_out_stage1[92]), .inData_93(wire_switch_out_stage1[93]), .inData_94(wire_switch_out_stage1[94]), .inData_95(wire_switch_out_stage1[95]), .inData_96(wire_switch_out_stage1[96]), .inData_97(wire_switch_out_stage1[97]), .inData_98(wire_switch_out_stage1[98]), .inData_99(wire_switch_out_stage1[99]), .inData_100(wire_switch_out_stage1[100]), .inData_101(wire_switch_out_stage1[101]), .inData_102(wire_switch_out_stage1[102]), .inData_103(wire_switch_out_stage1[103]), .inData_104(wire_switch_out_stage1[104]), .inData_105(wire_switch_out_stage1[105]), .inData_106(wire_switch_out_stage1[106]), .inData_107(wire_switch_out_stage1[107]), .inData_108(wire_switch_out_stage1[108]), .inData_109(wire_switch_out_stage1[109]), .inData_110(wire_switch_out_stage1[110]), .inData_111(wire_switch_out_stage1[111]), .inData_112(wire_switch_out_stage1[112]), .inData_113(wire_switch_out_stage1[113]), .inData_114(wire_switch_out_stage1[114]), .inData_115(wire_switch_out_stage1[115]), .inData_116(wire_switch_out_stage1[116]), .inData_117(wire_switch_out_stage1[117]), .inData_118(wire_switch_out_stage1[118]), .inData_119(wire_switch_out_stage1[119]), .inData_120(wire_switch_out_stage1[120]), .inData_121(wire_switch_out_stage1[121]), .inData_122(wire_switch_out_stage1[122]), .inData_123(wire_switch_out_stage1[123]), .inData_124(wire_switch_out_stage1[124]), .inData_125(wire_switch_out_stage1[125]), .inData_126(wire_switch_out_stage1[126]), .inData_127(wire_switch_out_stage1[127]), .inData_128(wire_switch_out_stage1[128]), .inData_129(wire_switch_out_stage1[129]), .inData_130(wire_switch_out_stage1[130]), .inData_131(wire_switch_out_stage1[131]), .inData_132(wire_switch_out_stage1[132]), .inData_133(wire_switch_out_stage1[133]), .inData_134(wire_switch_out_stage1[134]), .inData_135(wire_switch_out_stage1[135]), .inData_136(wire_switch_out_stage1[136]), .inData_137(wire_switch_out_stage1[137]), .inData_138(wire_switch_out_stage1[138]), .inData_139(wire_switch_out_stage1[139]), .inData_140(wire_switch_out_stage1[140]), .inData_141(wire_switch_out_stage1[141]), .inData_142(wire_switch_out_stage1[142]), .inData_143(wire_switch_out_stage1[143]), .inData_144(wire_switch_out_stage1[144]), .inData_145(wire_switch_out_stage1[145]), .inData_146(wire_switch_out_stage1[146]), .inData_147(wire_switch_out_stage1[147]), .inData_148(wire_switch_out_stage1[148]), .inData_149(wire_switch_out_stage1[149]), .inData_150(wire_switch_out_stage1[150]), .inData_151(wire_switch_out_stage1[151]), .inData_152(wire_switch_out_stage1[152]), .inData_153(wire_switch_out_stage1[153]), .inData_154(wire_switch_out_stage1[154]), .inData_155(wire_switch_out_stage1[155]), .inData_156(wire_switch_out_stage1[156]), .inData_157(wire_switch_out_stage1[157]), .inData_158(wire_switch_out_stage1[158]), .inData_159(wire_switch_out_stage1[159]), .inData_160(wire_switch_out_stage1[160]), .inData_161(wire_switch_out_stage1[161]), .inData_162(wire_switch_out_stage1[162]), .inData_163(wire_switch_out_stage1[163]), .inData_164(wire_switch_out_stage1[164]), .inData_165(wire_switch_out_stage1[165]), .inData_166(wire_switch_out_stage1[166]), .inData_167(wire_switch_out_stage1[167]), .inData_168(wire_switch_out_stage1[168]), .inData_169(wire_switch_out_stage1[169]), .inData_170(wire_switch_out_stage1[170]), .inData_171(wire_switch_out_stage1[171]), .inData_172(wire_switch_out_stage1[172]), .inData_173(wire_switch_out_stage1[173]), .inData_174(wire_switch_out_stage1[174]), .inData_175(wire_switch_out_stage1[175]), .inData_176(wire_switch_out_stage1[176]), .inData_177(wire_switch_out_stage1[177]), .inData_178(wire_switch_out_stage1[178]), .inData_179(wire_switch_out_stage1[179]), .inData_180(wire_switch_out_stage1[180]), .inData_181(wire_switch_out_stage1[181]), .inData_182(wire_switch_out_stage1[182]), .inData_183(wire_switch_out_stage1[183]), .inData_184(wire_switch_out_stage1[184]), .inData_185(wire_switch_out_stage1[185]), .inData_186(wire_switch_out_stage1[186]), .inData_187(wire_switch_out_stage1[187]), .inData_188(wire_switch_out_stage1[188]), .inData_189(wire_switch_out_stage1[189]), .inData_190(wire_switch_out_stage1[190]), .inData_191(wire_switch_out_stage1[191]), .inData_192(wire_switch_out_stage1[192]), .inData_193(wire_switch_out_stage1[193]), .inData_194(wire_switch_out_stage1[194]), .inData_195(wire_switch_out_stage1[195]), .inData_196(wire_switch_out_stage1[196]), .inData_197(wire_switch_out_stage1[197]), .inData_198(wire_switch_out_stage1[198]), .inData_199(wire_switch_out_stage1[199]), .inData_200(wire_switch_out_stage1[200]), .inData_201(wire_switch_out_stage1[201]), .inData_202(wire_switch_out_stage1[202]), .inData_203(wire_switch_out_stage1[203]), .inData_204(wire_switch_out_stage1[204]), .inData_205(wire_switch_out_stage1[205]), .inData_206(wire_switch_out_stage1[206]), .inData_207(wire_switch_out_stage1[207]), .inData_208(wire_switch_out_stage1[208]), .inData_209(wire_switch_out_stage1[209]), .inData_210(wire_switch_out_stage1[210]), .inData_211(wire_switch_out_stage1[211]), .inData_212(wire_switch_out_stage1[212]), .inData_213(wire_switch_out_stage1[213]), .inData_214(wire_switch_out_stage1[214]), .inData_215(wire_switch_out_stage1[215]), .inData_216(wire_switch_out_stage1[216]), .inData_217(wire_switch_out_stage1[217]), .inData_218(wire_switch_out_stage1[218]), .inData_219(wire_switch_out_stage1[219]), .inData_220(wire_switch_out_stage1[220]), .inData_221(wire_switch_out_stage1[221]), .inData_222(wire_switch_out_stage1[222]), .inData_223(wire_switch_out_stage1[223]), .inData_224(wire_switch_out_stage1[224]), .inData_225(wire_switch_out_stage1[225]), .inData_226(wire_switch_out_stage1[226]), .inData_227(wire_switch_out_stage1[227]), .inData_228(wire_switch_out_stage1[228]), .inData_229(wire_switch_out_stage1[229]), .inData_230(wire_switch_out_stage1[230]), .inData_231(wire_switch_out_stage1[231]), .inData_232(wire_switch_out_stage1[232]), .inData_233(wire_switch_out_stage1[233]), .inData_234(wire_switch_out_stage1[234]), .inData_235(wire_switch_out_stage1[235]), .inData_236(wire_switch_out_stage1[236]), .inData_237(wire_switch_out_stage1[237]), .inData_238(wire_switch_out_stage1[238]), .inData_239(wire_switch_out_stage1[239]), .inData_240(wire_switch_out_stage1[240]), .inData_241(wire_switch_out_stage1[241]), .inData_242(wire_switch_out_stage1[242]), .inData_243(wire_switch_out_stage1[243]), .inData_244(wire_switch_out_stage1[244]), .inData_245(wire_switch_out_stage1[245]), .inData_246(wire_switch_out_stage1[246]), .inData_247(wire_switch_out_stage1[247]), .inData_248(wire_switch_out_stage1[248]), .inData_249(wire_switch_out_stage1[249]), .inData_250(wire_switch_out_stage1[250]), .inData_251(wire_switch_out_stage1[251]), .inData_252(wire_switch_out_stage1[252]), .inData_253(wire_switch_out_stage1[253]), .inData_254(wire_switch_out_stage1[254]), .inData_255(wire_switch_out_stage1[255]), 
        .outData_0(wire_switch_in_stage0[0]), .outData_1(wire_switch_in_stage0[1]), .outData_2(wire_switch_in_stage0[2]), .outData_3(wire_switch_in_stage0[3]), .outData_4(wire_switch_in_stage0[4]), .outData_5(wire_switch_in_stage0[5]), .outData_6(wire_switch_in_stage0[6]), .outData_7(wire_switch_in_stage0[7]), .outData_8(wire_switch_in_stage0[8]), .outData_9(wire_switch_in_stage0[9]), .outData_10(wire_switch_in_stage0[10]), .outData_11(wire_switch_in_stage0[11]), .outData_12(wire_switch_in_stage0[12]), .outData_13(wire_switch_in_stage0[13]), .outData_14(wire_switch_in_stage0[14]), .outData_15(wire_switch_in_stage0[15]), .outData_16(wire_switch_in_stage0[16]), .outData_17(wire_switch_in_stage0[17]), .outData_18(wire_switch_in_stage0[18]), .outData_19(wire_switch_in_stage0[19]), .outData_20(wire_switch_in_stage0[20]), .outData_21(wire_switch_in_stage0[21]), .outData_22(wire_switch_in_stage0[22]), .outData_23(wire_switch_in_stage0[23]), .outData_24(wire_switch_in_stage0[24]), .outData_25(wire_switch_in_stage0[25]), .outData_26(wire_switch_in_stage0[26]), .outData_27(wire_switch_in_stage0[27]), .outData_28(wire_switch_in_stage0[28]), .outData_29(wire_switch_in_stage0[29]), .outData_30(wire_switch_in_stage0[30]), .outData_31(wire_switch_in_stage0[31]), .outData_32(wire_switch_in_stage0[32]), .outData_33(wire_switch_in_stage0[33]), .outData_34(wire_switch_in_stage0[34]), .outData_35(wire_switch_in_stage0[35]), .outData_36(wire_switch_in_stage0[36]), .outData_37(wire_switch_in_stage0[37]), .outData_38(wire_switch_in_stage0[38]), .outData_39(wire_switch_in_stage0[39]), .outData_40(wire_switch_in_stage0[40]), .outData_41(wire_switch_in_stage0[41]), .outData_42(wire_switch_in_stage0[42]), .outData_43(wire_switch_in_stage0[43]), .outData_44(wire_switch_in_stage0[44]), .outData_45(wire_switch_in_stage0[45]), .outData_46(wire_switch_in_stage0[46]), .outData_47(wire_switch_in_stage0[47]), .outData_48(wire_switch_in_stage0[48]), .outData_49(wire_switch_in_stage0[49]), .outData_50(wire_switch_in_stage0[50]), .outData_51(wire_switch_in_stage0[51]), .outData_52(wire_switch_in_stage0[52]), .outData_53(wire_switch_in_stage0[53]), .outData_54(wire_switch_in_stage0[54]), .outData_55(wire_switch_in_stage0[55]), .outData_56(wire_switch_in_stage0[56]), .outData_57(wire_switch_in_stage0[57]), .outData_58(wire_switch_in_stage0[58]), .outData_59(wire_switch_in_stage0[59]), .outData_60(wire_switch_in_stage0[60]), .outData_61(wire_switch_in_stage0[61]), .outData_62(wire_switch_in_stage0[62]), .outData_63(wire_switch_in_stage0[63]), .outData_64(wire_switch_in_stage0[64]), .outData_65(wire_switch_in_stage0[65]), .outData_66(wire_switch_in_stage0[66]), .outData_67(wire_switch_in_stage0[67]), .outData_68(wire_switch_in_stage0[68]), .outData_69(wire_switch_in_stage0[69]), .outData_70(wire_switch_in_stage0[70]), .outData_71(wire_switch_in_stage0[71]), .outData_72(wire_switch_in_stage0[72]), .outData_73(wire_switch_in_stage0[73]), .outData_74(wire_switch_in_stage0[74]), .outData_75(wire_switch_in_stage0[75]), .outData_76(wire_switch_in_stage0[76]), .outData_77(wire_switch_in_stage0[77]), .outData_78(wire_switch_in_stage0[78]), .outData_79(wire_switch_in_stage0[79]), .outData_80(wire_switch_in_stage0[80]), .outData_81(wire_switch_in_stage0[81]), .outData_82(wire_switch_in_stage0[82]), .outData_83(wire_switch_in_stage0[83]), .outData_84(wire_switch_in_stage0[84]), .outData_85(wire_switch_in_stage0[85]), .outData_86(wire_switch_in_stage0[86]), .outData_87(wire_switch_in_stage0[87]), .outData_88(wire_switch_in_stage0[88]), .outData_89(wire_switch_in_stage0[89]), .outData_90(wire_switch_in_stage0[90]), .outData_91(wire_switch_in_stage0[91]), .outData_92(wire_switch_in_stage0[92]), .outData_93(wire_switch_in_stage0[93]), .outData_94(wire_switch_in_stage0[94]), .outData_95(wire_switch_in_stage0[95]), .outData_96(wire_switch_in_stage0[96]), .outData_97(wire_switch_in_stage0[97]), .outData_98(wire_switch_in_stage0[98]), .outData_99(wire_switch_in_stage0[99]), .outData_100(wire_switch_in_stage0[100]), .outData_101(wire_switch_in_stage0[101]), .outData_102(wire_switch_in_stage0[102]), .outData_103(wire_switch_in_stage0[103]), .outData_104(wire_switch_in_stage0[104]), .outData_105(wire_switch_in_stage0[105]), .outData_106(wire_switch_in_stage0[106]), .outData_107(wire_switch_in_stage0[107]), .outData_108(wire_switch_in_stage0[108]), .outData_109(wire_switch_in_stage0[109]), .outData_110(wire_switch_in_stage0[110]), .outData_111(wire_switch_in_stage0[111]), .outData_112(wire_switch_in_stage0[112]), .outData_113(wire_switch_in_stage0[113]), .outData_114(wire_switch_in_stage0[114]), .outData_115(wire_switch_in_stage0[115]), .outData_116(wire_switch_in_stage0[116]), .outData_117(wire_switch_in_stage0[117]), .outData_118(wire_switch_in_stage0[118]), .outData_119(wire_switch_in_stage0[119]), .outData_120(wire_switch_in_stage0[120]), .outData_121(wire_switch_in_stage0[121]), .outData_122(wire_switch_in_stage0[122]), .outData_123(wire_switch_in_stage0[123]), .outData_124(wire_switch_in_stage0[124]), .outData_125(wire_switch_in_stage0[125]), .outData_126(wire_switch_in_stage0[126]), .outData_127(wire_switch_in_stage0[127]), .outData_128(wire_switch_in_stage0[128]), .outData_129(wire_switch_in_stage0[129]), .outData_130(wire_switch_in_stage0[130]), .outData_131(wire_switch_in_stage0[131]), .outData_132(wire_switch_in_stage0[132]), .outData_133(wire_switch_in_stage0[133]), .outData_134(wire_switch_in_stage0[134]), .outData_135(wire_switch_in_stage0[135]), .outData_136(wire_switch_in_stage0[136]), .outData_137(wire_switch_in_stage0[137]), .outData_138(wire_switch_in_stage0[138]), .outData_139(wire_switch_in_stage0[139]), .outData_140(wire_switch_in_stage0[140]), .outData_141(wire_switch_in_stage0[141]), .outData_142(wire_switch_in_stage0[142]), .outData_143(wire_switch_in_stage0[143]), .outData_144(wire_switch_in_stage0[144]), .outData_145(wire_switch_in_stage0[145]), .outData_146(wire_switch_in_stage0[146]), .outData_147(wire_switch_in_stage0[147]), .outData_148(wire_switch_in_stage0[148]), .outData_149(wire_switch_in_stage0[149]), .outData_150(wire_switch_in_stage0[150]), .outData_151(wire_switch_in_stage0[151]), .outData_152(wire_switch_in_stage0[152]), .outData_153(wire_switch_in_stage0[153]), .outData_154(wire_switch_in_stage0[154]), .outData_155(wire_switch_in_stage0[155]), .outData_156(wire_switch_in_stage0[156]), .outData_157(wire_switch_in_stage0[157]), .outData_158(wire_switch_in_stage0[158]), .outData_159(wire_switch_in_stage0[159]), .outData_160(wire_switch_in_stage0[160]), .outData_161(wire_switch_in_stage0[161]), .outData_162(wire_switch_in_stage0[162]), .outData_163(wire_switch_in_stage0[163]), .outData_164(wire_switch_in_stage0[164]), .outData_165(wire_switch_in_stage0[165]), .outData_166(wire_switch_in_stage0[166]), .outData_167(wire_switch_in_stage0[167]), .outData_168(wire_switch_in_stage0[168]), .outData_169(wire_switch_in_stage0[169]), .outData_170(wire_switch_in_stage0[170]), .outData_171(wire_switch_in_stage0[171]), .outData_172(wire_switch_in_stage0[172]), .outData_173(wire_switch_in_stage0[173]), .outData_174(wire_switch_in_stage0[174]), .outData_175(wire_switch_in_stage0[175]), .outData_176(wire_switch_in_stage0[176]), .outData_177(wire_switch_in_stage0[177]), .outData_178(wire_switch_in_stage0[178]), .outData_179(wire_switch_in_stage0[179]), .outData_180(wire_switch_in_stage0[180]), .outData_181(wire_switch_in_stage0[181]), .outData_182(wire_switch_in_stage0[182]), .outData_183(wire_switch_in_stage0[183]), .outData_184(wire_switch_in_stage0[184]), .outData_185(wire_switch_in_stage0[185]), .outData_186(wire_switch_in_stage0[186]), .outData_187(wire_switch_in_stage0[187]), .outData_188(wire_switch_in_stage0[188]), .outData_189(wire_switch_in_stage0[189]), .outData_190(wire_switch_in_stage0[190]), .outData_191(wire_switch_in_stage0[191]), .outData_192(wire_switch_in_stage0[192]), .outData_193(wire_switch_in_stage0[193]), .outData_194(wire_switch_in_stage0[194]), .outData_195(wire_switch_in_stage0[195]), .outData_196(wire_switch_in_stage0[196]), .outData_197(wire_switch_in_stage0[197]), .outData_198(wire_switch_in_stage0[198]), .outData_199(wire_switch_in_stage0[199]), .outData_200(wire_switch_in_stage0[200]), .outData_201(wire_switch_in_stage0[201]), .outData_202(wire_switch_in_stage0[202]), .outData_203(wire_switch_in_stage0[203]), .outData_204(wire_switch_in_stage0[204]), .outData_205(wire_switch_in_stage0[205]), .outData_206(wire_switch_in_stage0[206]), .outData_207(wire_switch_in_stage0[207]), .outData_208(wire_switch_in_stage0[208]), .outData_209(wire_switch_in_stage0[209]), .outData_210(wire_switch_in_stage0[210]), .outData_211(wire_switch_in_stage0[211]), .outData_212(wire_switch_in_stage0[212]), .outData_213(wire_switch_in_stage0[213]), .outData_214(wire_switch_in_stage0[214]), .outData_215(wire_switch_in_stage0[215]), .outData_216(wire_switch_in_stage0[216]), .outData_217(wire_switch_in_stage0[217]), .outData_218(wire_switch_in_stage0[218]), .outData_219(wire_switch_in_stage0[219]), .outData_220(wire_switch_in_stage0[220]), .outData_221(wire_switch_in_stage0[221]), .outData_222(wire_switch_in_stage0[222]), .outData_223(wire_switch_in_stage0[223]), .outData_224(wire_switch_in_stage0[224]), .outData_225(wire_switch_in_stage0[225]), .outData_226(wire_switch_in_stage0[226]), .outData_227(wire_switch_in_stage0[227]), .outData_228(wire_switch_in_stage0[228]), .outData_229(wire_switch_in_stage0[229]), .outData_230(wire_switch_in_stage0[230]), .outData_231(wire_switch_in_stage0[231]), .outData_232(wire_switch_in_stage0[232]), .outData_233(wire_switch_in_stage0[233]), .outData_234(wire_switch_in_stage0[234]), .outData_235(wire_switch_in_stage0[235]), .outData_236(wire_switch_in_stage0[236]), .outData_237(wire_switch_in_stage0[237]), .outData_238(wire_switch_in_stage0[238]), .outData_239(wire_switch_in_stage0[239]), .outData_240(wire_switch_in_stage0[240]), .outData_241(wire_switch_in_stage0[241]), .outData_242(wire_switch_in_stage0[242]), .outData_243(wire_switch_in_stage0[243]), .outData_244(wire_switch_in_stage0[244]), .outData_245(wire_switch_in_stage0[245]), .outData_246(wire_switch_in_stage0[246]), .outData_247(wire_switch_in_stage0[247]), .outData_248(wire_switch_in_stage0[248]), .outData_249(wire_switch_in_stage0[249]), .outData_250(wire_switch_in_stage0[250]), .outData_251(wire_switch_in_stage0[251]), .outData_252(wire_switch_in_stage0[252]), .outData_253(wire_switch_in_stage0[253]), .outData_254(wire_switch_in_stage0[254]), .outData_255(wire_switch_in_stage0[255]), 
        .in_start(in_start_stage0), .out_start(con_in_start_stage0), .clk(clk), .rst(rst)); 

  
  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[0] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[1] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[2] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[3] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[4] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[5] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[6] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[7] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[8] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[9] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[10] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[11] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[12] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[13] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[14] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[15] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[16] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[17] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[18] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[19] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[20] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[21] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[22] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[23] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[24] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[25] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[26] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[27] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[28] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[29] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[30] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[31] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[32] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[33] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[34] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[35] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[36] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[37] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[38] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[39] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[40] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[41] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[42] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[43] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[44] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[45] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[46] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[47] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[48] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[49] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[50] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[51] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[52] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[53] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[54] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[55] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[56] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[57] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[58] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[59] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[60] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[61] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[62] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[63] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[64] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[65] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[66] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[67] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[68] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[69] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[70] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[71] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[72] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[73] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[74] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[75] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[76] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[77] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[78] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[79] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[80] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[81] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[82] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[83] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[84] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[85] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[86] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[87] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[88] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[89] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[90] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[91] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[92] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[93] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[94] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[95] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[96] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[97] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[98] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[99] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[100] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[101] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[102] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[103] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[104] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[105] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[106] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[107] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[108] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[109] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[110] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[111] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[112] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[113] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[114] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[115] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[116] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[117] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[118] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[119] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[120] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[121] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[122] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[123] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[124] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[125] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[126] <= counter_w[7]; 
  end                            

  always@(posedge clk)             
  begin                            
    wire_ctrl_stage0[127] <= counter_w[7]; 
  end                            

  
  assign in_start_stage7 = in_start;    
  assign outData_0 = wireOut[0];    
  assign outData_1 = wireOut[1];    
  assign outData_2 = wireOut[2];    
  assign outData_3 = wireOut[3];    
  assign outData_4 = wireOut[4];    
  assign outData_5 = wireOut[5];    
  assign outData_6 = wireOut[6];    
  assign outData_7 = wireOut[7];    
  assign outData_8 = wireOut[8];    
  assign outData_9 = wireOut[9];    
  assign outData_10 = wireOut[10];    
  assign outData_11 = wireOut[11];    
  assign outData_12 = wireOut[12];    
  assign outData_13 = wireOut[13];    
  assign outData_14 = wireOut[14];    
  assign outData_15 = wireOut[15];    
  assign outData_16 = wireOut[16];    
  assign outData_17 = wireOut[17];    
  assign outData_18 = wireOut[18];    
  assign outData_19 = wireOut[19];    
  assign outData_20 = wireOut[20];    
  assign outData_21 = wireOut[21];    
  assign outData_22 = wireOut[22];    
  assign outData_23 = wireOut[23];    
  assign outData_24 = wireOut[24];    
  assign outData_25 = wireOut[25];    
  assign outData_26 = wireOut[26];    
  assign outData_27 = wireOut[27];    
  assign outData_28 = wireOut[28];    
  assign outData_29 = wireOut[29];    
  assign outData_30 = wireOut[30];    
  assign outData_31 = wireOut[31];    
  assign outData_32 = wireOut[32];    
  assign outData_33 = wireOut[33];    
  assign outData_34 = wireOut[34];    
  assign outData_35 = wireOut[35];    
  assign outData_36 = wireOut[36];    
  assign outData_37 = wireOut[37];    
  assign outData_38 = wireOut[38];    
  assign outData_39 = wireOut[39];    
  assign outData_40 = wireOut[40];    
  assign outData_41 = wireOut[41];    
  assign outData_42 = wireOut[42];    
  assign outData_43 = wireOut[43];    
  assign outData_44 = wireOut[44];    
  assign outData_45 = wireOut[45];    
  assign outData_46 = wireOut[46];    
  assign outData_47 = wireOut[47];    
  assign outData_48 = wireOut[48];    
  assign outData_49 = wireOut[49];    
  assign outData_50 = wireOut[50];    
  assign outData_51 = wireOut[51];    
  assign outData_52 = wireOut[52];    
  assign outData_53 = wireOut[53];    
  assign outData_54 = wireOut[54];    
  assign outData_55 = wireOut[55];    
  assign outData_56 = wireOut[56];    
  assign outData_57 = wireOut[57];    
  assign outData_58 = wireOut[58];    
  assign outData_59 = wireOut[59];    
  assign outData_60 = wireOut[60];    
  assign outData_61 = wireOut[61];    
  assign outData_62 = wireOut[62];    
  assign outData_63 = wireOut[63];    
  assign outData_64 = wireOut[64];    
  assign outData_65 = wireOut[65];    
  assign outData_66 = wireOut[66];    
  assign outData_67 = wireOut[67];    
  assign outData_68 = wireOut[68];    
  assign outData_69 = wireOut[69];    
  assign outData_70 = wireOut[70];    
  assign outData_71 = wireOut[71];    
  assign outData_72 = wireOut[72];    
  assign outData_73 = wireOut[73];    
  assign outData_74 = wireOut[74];    
  assign outData_75 = wireOut[75];    
  assign outData_76 = wireOut[76];    
  assign outData_77 = wireOut[77];    
  assign outData_78 = wireOut[78];    
  assign outData_79 = wireOut[79];    
  assign outData_80 = wireOut[80];    
  assign outData_81 = wireOut[81];    
  assign outData_82 = wireOut[82];    
  assign outData_83 = wireOut[83];    
  assign outData_84 = wireOut[84];    
  assign outData_85 = wireOut[85];    
  assign outData_86 = wireOut[86];    
  assign outData_87 = wireOut[87];    
  assign outData_88 = wireOut[88];    
  assign outData_89 = wireOut[89];    
  assign outData_90 = wireOut[90];    
  assign outData_91 = wireOut[91];    
  assign outData_92 = wireOut[92];    
  assign outData_93 = wireOut[93];    
  assign outData_94 = wireOut[94];    
  assign outData_95 = wireOut[95];    
  assign outData_96 = wireOut[96];    
  assign outData_97 = wireOut[97];    
  assign outData_98 = wireOut[98];    
  assign outData_99 = wireOut[99];    
  assign outData_100 = wireOut[100];    
  assign outData_101 = wireOut[101];    
  assign outData_102 = wireOut[102];    
  assign outData_103 = wireOut[103];    
  assign outData_104 = wireOut[104];    
  assign outData_105 = wireOut[105];    
  assign outData_106 = wireOut[106];    
  assign outData_107 = wireOut[107];    
  assign outData_108 = wireOut[108];    
  assign outData_109 = wireOut[109];    
  assign outData_110 = wireOut[110];    
  assign outData_111 = wireOut[111];    
  assign outData_112 = wireOut[112];    
  assign outData_113 = wireOut[113];    
  assign outData_114 = wireOut[114];    
  assign outData_115 = wireOut[115];    
  assign outData_116 = wireOut[116];    
  assign outData_117 = wireOut[117];    
  assign outData_118 = wireOut[118];    
  assign outData_119 = wireOut[119];    
  assign outData_120 = wireOut[120];    
  assign outData_121 = wireOut[121];    
  assign outData_122 = wireOut[122];    
  assign outData_123 = wireOut[123];    
  assign outData_124 = wireOut[124];    
  assign outData_125 = wireOut[125];    
  assign outData_126 = wireOut[126];    
  assign outData_127 = wireOut[127];    
  assign outData_128 = wireOut[128];    
  assign outData_129 = wireOut[129];    
  assign outData_130 = wireOut[130];    
  assign outData_131 = wireOut[131];    
  assign outData_132 = wireOut[132];    
  assign outData_133 = wireOut[133];    
  assign outData_134 = wireOut[134];    
  assign outData_135 = wireOut[135];    
  assign outData_136 = wireOut[136];    
  assign outData_137 = wireOut[137];    
  assign outData_138 = wireOut[138];    
  assign outData_139 = wireOut[139];    
  assign outData_140 = wireOut[140];    
  assign outData_141 = wireOut[141];    
  assign outData_142 = wireOut[142];    
  assign outData_143 = wireOut[143];    
  assign outData_144 = wireOut[144];    
  assign outData_145 = wireOut[145];    
  assign outData_146 = wireOut[146];    
  assign outData_147 = wireOut[147];    
  assign outData_148 = wireOut[148];    
  assign outData_149 = wireOut[149];    
  assign outData_150 = wireOut[150];    
  assign outData_151 = wireOut[151];    
  assign outData_152 = wireOut[152];    
  assign outData_153 = wireOut[153];    
  assign outData_154 = wireOut[154];    
  assign outData_155 = wireOut[155];    
  assign outData_156 = wireOut[156];    
  assign outData_157 = wireOut[157];    
  assign outData_158 = wireOut[158];    
  assign outData_159 = wireOut[159];    
  assign outData_160 = wireOut[160];    
  assign outData_161 = wireOut[161];    
  assign outData_162 = wireOut[162];    
  assign outData_163 = wireOut[163];    
  assign outData_164 = wireOut[164];    
  assign outData_165 = wireOut[165];    
  assign outData_166 = wireOut[166];    
  assign outData_167 = wireOut[167];    
  assign outData_168 = wireOut[168];    
  assign outData_169 = wireOut[169];    
  assign outData_170 = wireOut[170];    
  assign outData_171 = wireOut[171];    
  assign outData_172 = wireOut[172];    
  assign outData_173 = wireOut[173];    
  assign outData_174 = wireOut[174];    
  assign outData_175 = wireOut[175];    
  assign outData_176 = wireOut[176];    
  assign outData_177 = wireOut[177];    
  assign outData_178 = wireOut[178];    
  assign outData_179 = wireOut[179];    
  assign outData_180 = wireOut[180];    
  assign outData_181 = wireOut[181];    
  assign outData_182 = wireOut[182];    
  assign outData_183 = wireOut[183];    
  assign outData_184 = wireOut[184];    
  assign outData_185 = wireOut[185];    
  assign outData_186 = wireOut[186];    
  assign outData_187 = wireOut[187];    
  assign outData_188 = wireOut[188];    
  assign outData_189 = wireOut[189];    
  assign outData_190 = wireOut[190];    
  assign outData_191 = wireOut[191];    
  assign outData_192 = wireOut[192];    
  assign outData_193 = wireOut[193];    
  assign outData_194 = wireOut[194];    
  assign outData_195 = wireOut[195];    
  assign outData_196 = wireOut[196];    
  assign outData_197 = wireOut[197];    
  assign outData_198 = wireOut[198];    
  assign outData_199 = wireOut[199];    
  assign outData_200 = wireOut[200];    
  assign outData_201 = wireOut[201];    
  assign outData_202 = wireOut[202];    
  assign outData_203 = wireOut[203];    
  assign outData_204 = wireOut[204];    
  assign outData_205 = wireOut[205];    
  assign outData_206 = wireOut[206];    
  assign outData_207 = wireOut[207];    
  assign outData_208 = wireOut[208];    
  assign outData_209 = wireOut[209];    
  assign outData_210 = wireOut[210];    
  assign outData_211 = wireOut[211];    
  assign outData_212 = wireOut[212];    
  assign outData_213 = wireOut[213];    
  assign outData_214 = wireOut[214];    
  assign outData_215 = wireOut[215];    
  assign outData_216 = wireOut[216];    
  assign outData_217 = wireOut[217];    
  assign outData_218 = wireOut[218];    
  assign outData_219 = wireOut[219];    
  assign outData_220 = wireOut[220];    
  assign outData_221 = wireOut[221];    
  assign outData_222 = wireOut[222];    
  assign outData_223 = wireOut[223];    
  assign outData_224 = wireOut[224];    
  assign outData_225 = wireOut[225];    
  assign outData_226 = wireOut[226];    
  assign outData_227 = wireOut[227];    
  assign outData_228 = wireOut[228];    
  assign outData_229 = wireOut[229];    
  assign outData_230 = wireOut[230];    
  assign outData_231 = wireOut[231];    
  assign outData_232 = wireOut[232];    
  assign outData_233 = wireOut[233];    
  assign outData_234 = wireOut[234];    
  assign outData_235 = wireOut[235];    
  assign outData_236 = wireOut[236];    
  assign outData_237 = wireOut[237];    
  assign outData_238 = wireOut[238];    
  assign outData_239 = wireOut[239];    
  assign outData_240 = wireOut[240];    
  assign outData_241 = wireOut[241];    
  assign outData_242 = wireOut[242];    
  assign outData_243 = wireOut[243];    
  assign outData_244 = wireOut[244];    
  assign outData_245 = wireOut[245];    
  assign outData_246 = wireOut[246];    
  assign outData_247 = wireOut[247];    
  assign outData_248 = wireOut[248];    
  assign outData_249 = wireOut[249];    
  assign outData_250 = wireOut[250];    
  assign outData_251 = wireOut[251];    
  assign outData_252 = wireOut[252];    
  assign outData_253 = wireOut[253];    
  assign outData_254 = wireOut[254];    
  assign outData_255 = wireOut[255];    
  assign out_start = out_start_w;    
  
endmodule                        


module  mem_addr_gen_dp256_mem0_per0(
counter_in,                              
clk,                             
rst,                             
addr_out                            
);                               
  input clk, rst;                           
  input [7:0] counter_in;      
  output [7:0] addr_out;      

  wire [7:0] addr_a0;      
  assign addr_out[7:0] = addr_a0[7:0];   
  
  assign addr_a0 = counter_in[7:0]; 
  
endmodule                        


module  mem_addr_ctrl_dp256_per0(
in_start,                          
counter_in,                         
wen_out,                         
out_start,                         
mem_addr_out_0,                         
mem_addr_out_1,                         
mem_addr_out_2,                         
mem_addr_out_3,                         
mem_addr_out_4,                         
mem_addr_out_5,                         
mem_addr_out_6,                         
mem_addr_out_7,                         
mem_addr_out_8,                         
mem_addr_out_9,                         
mem_addr_out_10,                         
mem_addr_out_11,                         
mem_addr_out_12,                         
mem_addr_out_13,                         
mem_addr_out_14,                         
mem_addr_out_15,                         
mem_addr_out_16,                         
mem_addr_out_17,                         
mem_addr_out_18,                         
mem_addr_out_19,                         
mem_addr_out_20,                         
mem_addr_out_21,                         
mem_addr_out_22,                         
mem_addr_out_23,                         
mem_addr_out_24,                         
mem_addr_out_25,                         
mem_addr_out_26,                         
mem_addr_out_27,                         
mem_addr_out_28,                         
mem_addr_out_29,                         
mem_addr_out_30,                         
mem_addr_out_31,                         
mem_addr_out_32,                         
mem_addr_out_33,                         
mem_addr_out_34,                         
mem_addr_out_35,                         
mem_addr_out_36,                         
mem_addr_out_37,                         
mem_addr_out_38,                         
mem_addr_out_39,                         
mem_addr_out_40,                         
mem_addr_out_41,                         
mem_addr_out_42,                         
mem_addr_out_43,                         
mem_addr_out_44,                         
mem_addr_out_45,                         
mem_addr_out_46,                         
mem_addr_out_47,                         
mem_addr_out_48,                         
mem_addr_out_49,                         
mem_addr_out_50,                         
mem_addr_out_51,                         
mem_addr_out_52,                         
mem_addr_out_53,                         
mem_addr_out_54,                         
mem_addr_out_55,                         
mem_addr_out_56,                         
mem_addr_out_57,                         
mem_addr_out_58,                         
mem_addr_out_59,                         
mem_addr_out_60,                         
mem_addr_out_61,                         
mem_addr_out_62,                         
mem_addr_out_63,                         
mem_addr_out_64,                         
mem_addr_out_65,                         
mem_addr_out_66,                         
mem_addr_out_67,                         
mem_addr_out_68,                         
mem_addr_out_69,                         
mem_addr_out_70,                         
mem_addr_out_71,                         
mem_addr_out_72,                         
mem_addr_out_73,                         
mem_addr_out_74,                         
mem_addr_out_75,                         
mem_addr_out_76,                         
mem_addr_out_77,                         
mem_addr_out_78,                         
mem_addr_out_79,                         
mem_addr_out_80,                         
mem_addr_out_81,                         
mem_addr_out_82,                         
mem_addr_out_83,                         
mem_addr_out_84,                         
mem_addr_out_85,                         
mem_addr_out_86,                         
mem_addr_out_87,                         
mem_addr_out_88,                         
mem_addr_out_89,                         
mem_addr_out_90,                         
mem_addr_out_91,                         
mem_addr_out_92,                         
mem_addr_out_93,                         
mem_addr_out_94,                         
mem_addr_out_95,                         
mem_addr_out_96,                         
mem_addr_out_97,                         
mem_addr_out_98,                         
mem_addr_out_99,                         
mem_addr_out_100,                         
mem_addr_out_101,                         
mem_addr_out_102,                         
mem_addr_out_103,                         
mem_addr_out_104,                         
mem_addr_out_105,                         
mem_addr_out_106,                         
mem_addr_out_107,                         
mem_addr_out_108,                         
mem_addr_out_109,                         
mem_addr_out_110,                         
mem_addr_out_111,                         
mem_addr_out_112,                         
mem_addr_out_113,                         
mem_addr_out_114,                         
mem_addr_out_115,                         
mem_addr_out_116,                         
mem_addr_out_117,                         
mem_addr_out_118,                         
mem_addr_out_119,                         
mem_addr_out_120,                         
mem_addr_out_121,                         
mem_addr_out_122,                         
mem_addr_out_123,                         
mem_addr_out_124,                         
mem_addr_out_125,                         
mem_addr_out_126,                         
mem_addr_out_127,                         
mem_addr_out_128,                         
mem_addr_out_129,                         
mem_addr_out_130,                         
mem_addr_out_131,                         
mem_addr_out_132,                         
mem_addr_out_133,                         
mem_addr_out_134,                         
mem_addr_out_135,                         
mem_addr_out_136,                         
mem_addr_out_137,                         
mem_addr_out_138,                         
mem_addr_out_139,                         
mem_addr_out_140,                         
mem_addr_out_141,                         
mem_addr_out_142,                         
mem_addr_out_143,                         
mem_addr_out_144,                         
mem_addr_out_145,                         
mem_addr_out_146,                         
mem_addr_out_147,                         
mem_addr_out_148,                         
mem_addr_out_149,                         
mem_addr_out_150,                         
mem_addr_out_151,                         
mem_addr_out_152,                         
mem_addr_out_153,                         
mem_addr_out_154,                         
mem_addr_out_155,                         
mem_addr_out_156,                         
mem_addr_out_157,                         
mem_addr_out_158,                         
mem_addr_out_159,                         
mem_addr_out_160,                         
mem_addr_out_161,                         
mem_addr_out_162,                         
mem_addr_out_163,                         
mem_addr_out_164,                         
mem_addr_out_165,                         
mem_addr_out_166,                         
mem_addr_out_167,                         
mem_addr_out_168,                         
mem_addr_out_169,                         
mem_addr_out_170,                         
mem_addr_out_171,                         
mem_addr_out_172,                         
mem_addr_out_173,                         
mem_addr_out_174,                         
mem_addr_out_175,                         
mem_addr_out_176,                         
mem_addr_out_177,                         
mem_addr_out_178,                         
mem_addr_out_179,                         
mem_addr_out_180,                         
mem_addr_out_181,                         
mem_addr_out_182,                         
mem_addr_out_183,                         
mem_addr_out_184,                         
mem_addr_out_185,                         
mem_addr_out_186,                         
mem_addr_out_187,                         
mem_addr_out_188,                         
mem_addr_out_189,                         
mem_addr_out_190,                         
mem_addr_out_191,                         
mem_addr_out_192,                         
mem_addr_out_193,                         
mem_addr_out_194,                         
mem_addr_out_195,                         
mem_addr_out_196,                         
mem_addr_out_197,                         
mem_addr_out_198,                         
mem_addr_out_199,                         
mem_addr_out_200,                         
mem_addr_out_201,                         
mem_addr_out_202,                         
mem_addr_out_203,                         
mem_addr_out_204,                         
mem_addr_out_205,                         
mem_addr_out_206,                         
mem_addr_out_207,                         
mem_addr_out_208,                         
mem_addr_out_209,                         
mem_addr_out_210,                         
mem_addr_out_211,                         
mem_addr_out_212,                         
mem_addr_out_213,                         
mem_addr_out_214,                         
mem_addr_out_215,                         
mem_addr_out_216,                         
mem_addr_out_217,                         
mem_addr_out_218,                         
mem_addr_out_219,                         
mem_addr_out_220,                         
mem_addr_out_221,                         
mem_addr_out_222,                         
mem_addr_out_223,                         
mem_addr_out_224,                         
mem_addr_out_225,                         
mem_addr_out_226,                         
mem_addr_out_227,                         
mem_addr_out_228,                         
mem_addr_out_229,                         
mem_addr_out_230,                         
mem_addr_out_231,                         
mem_addr_out_232,                         
mem_addr_out_233,                         
mem_addr_out_234,                         
mem_addr_out_235,                         
mem_addr_out_236,                         
mem_addr_out_237,                         
mem_addr_out_238,                         
mem_addr_out_239,                         
mem_addr_out_240,                         
mem_addr_out_241,                         
mem_addr_out_242,                         
mem_addr_out_243,                         
mem_addr_out_244,                         
mem_addr_out_245,                         
mem_addr_out_246,                         
mem_addr_out_247,                         
mem_addr_out_248,                         
mem_addr_out_249,                         
mem_addr_out_250,                         
mem_addr_out_251,                         
mem_addr_out_252,                         
mem_addr_out_253,                         
mem_addr_out_254,                         
mem_addr_out_255,                         
clk,                             
rst                              
);                               
  input in_start, clk, rst;                   
  input [7:0] counter_in; 
  output [7:0] mem_addr_out_0;            
  output [7:0] mem_addr_out_1;            
  output [7:0] mem_addr_out_2;            
  output [7:0] mem_addr_out_3;            
  output [7:0] mem_addr_out_4;            
  output [7:0] mem_addr_out_5;            
  output [7:0] mem_addr_out_6;            
  output [7:0] mem_addr_out_7;            
  output [7:0] mem_addr_out_8;            
  output [7:0] mem_addr_out_9;            
  output [7:0] mem_addr_out_10;            
  output [7:0] mem_addr_out_11;            
  output [7:0] mem_addr_out_12;            
  output [7:0] mem_addr_out_13;            
  output [7:0] mem_addr_out_14;            
  output [7:0] mem_addr_out_15;            
  output [7:0] mem_addr_out_16;            
  output [7:0] mem_addr_out_17;            
  output [7:0] mem_addr_out_18;            
  output [7:0] mem_addr_out_19;            
  output [7:0] mem_addr_out_20;            
  output [7:0] mem_addr_out_21;            
  output [7:0] mem_addr_out_22;            
  output [7:0] mem_addr_out_23;            
  output [7:0] mem_addr_out_24;            
  output [7:0] mem_addr_out_25;            
  output [7:0] mem_addr_out_26;            
  output [7:0] mem_addr_out_27;            
  output [7:0] mem_addr_out_28;            
  output [7:0] mem_addr_out_29;            
  output [7:0] mem_addr_out_30;            
  output [7:0] mem_addr_out_31;            
  output [7:0] mem_addr_out_32;            
  output [7:0] mem_addr_out_33;            
  output [7:0] mem_addr_out_34;            
  output [7:0] mem_addr_out_35;            
  output [7:0] mem_addr_out_36;            
  output [7:0] mem_addr_out_37;            
  output [7:0] mem_addr_out_38;            
  output [7:0] mem_addr_out_39;            
  output [7:0] mem_addr_out_40;            
  output [7:0] mem_addr_out_41;            
  output [7:0] mem_addr_out_42;            
  output [7:0] mem_addr_out_43;            
  output [7:0] mem_addr_out_44;            
  output [7:0] mem_addr_out_45;            
  output [7:0] mem_addr_out_46;            
  output [7:0] mem_addr_out_47;            
  output [7:0] mem_addr_out_48;            
  output [7:0] mem_addr_out_49;            
  output [7:0] mem_addr_out_50;            
  output [7:0] mem_addr_out_51;            
  output [7:0] mem_addr_out_52;            
  output [7:0] mem_addr_out_53;            
  output [7:0] mem_addr_out_54;            
  output [7:0] mem_addr_out_55;            
  output [7:0] mem_addr_out_56;            
  output [7:0] mem_addr_out_57;            
  output [7:0] mem_addr_out_58;            
  output [7:0] mem_addr_out_59;            
  output [7:0] mem_addr_out_60;            
  output [7:0] mem_addr_out_61;            
  output [7:0] mem_addr_out_62;            
  output [7:0] mem_addr_out_63;            
  output [7:0] mem_addr_out_64;            
  output [7:0] mem_addr_out_65;            
  output [7:0] mem_addr_out_66;            
  output [7:0] mem_addr_out_67;            
  output [7:0] mem_addr_out_68;            
  output [7:0] mem_addr_out_69;            
  output [7:0] mem_addr_out_70;            
  output [7:0] mem_addr_out_71;            
  output [7:0] mem_addr_out_72;            
  output [7:0] mem_addr_out_73;            
  output [7:0] mem_addr_out_74;            
  output [7:0] mem_addr_out_75;            
  output [7:0] mem_addr_out_76;            
  output [7:0] mem_addr_out_77;            
  output [7:0] mem_addr_out_78;            
  output [7:0] mem_addr_out_79;            
  output [7:0] mem_addr_out_80;            
  output [7:0] mem_addr_out_81;            
  output [7:0] mem_addr_out_82;            
  output [7:0] mem_addr_out_83;            
  output [7:0] mem_addr_out_84;            
  output [7:0] mem_addr_out_85;            
  output [7:0] mem_addr_out_86;            
  output [7:0] mem_addr_out_87;            
  output [7:0] mem_addr_out_88;            
  output [7:0] mem_addr_out_89;            
  output [7:0] mem_addr_out_90;            
  output [7:0] mem_addr_out_91;            
  output [7:0] mem_addr_out_92;            
  output [7:0] mem_addr_out_93;            
  output [7:0] mem_addr_out_94;            
  output [7:0] mem_addr_out_95;            
  output [7:0] mem_addr_out_96;            
  output [7:0] mem_addr_out_97;            
  output [7:0] mem_addr_out_98;            
  output [7:0] mem_addr_out_99;            
  output [7:0] mem_addr_out_100;            
  output [7:0] mem_addr_out_101;            
  output [7:0] mem_addr_out_102;            
  output [7:0] mem_addr_out_103;            
  output [7:0] mem_addr_out_104;            
  output [7:0] mem_addr_out_105;            
  output [7:0] mem_addr_out_106;            
  output [7:0] mem_addr_out_107;            
  output [7:0] mem_addr_out_108;            
  output [7:0] mem_addr_out_109;            
  output [7:0] mem_addr_out_110;            
  output [7:0] mem_addr_out_111;            
  output [7:0] mem_addr_out_112;            
  output [7:0] mem_addr_out_113;            
  output [7:0] mem_addr_out_114;            
  output [7:0] mem_addr_out_115;            
  output [7:0] mem_addr_out_116;            
  output [7:0] mem_addr_out_117;            
  output [7:0] mem_addr_out_118;            
  output [7:0] mem_addr_out_119;            
  output [7:0] mem_addr_out_120;            
  output [7:0] mem_addr_out_121;            
  output [7:0] mem_addr_out_122;            
  output [7:0] mem_addr_out_123;            
  output [7:0] mem_addr_out_124;            
  output [7:0] mem_addr_out_125;            
  output [7:0] mem_addr_out_126;            
  output [7:0] mem_addr_out_127;            
  output [7:0] mem_addr_out_128;            
  output [7:0] mem_addr_out_129;            
  output [7:0] mem_addr_out_130;            
  output [7:0] mem_addr_out_131;            
  output [7:0] mem_addr_out_132;            
  output [7:0] mem_addr_out_133;            
  output [7:0] mem_addr_out_134;            
  output [7:0] mem_addr_out_135;            
  output [7:0] mem_addr_out_136;            
  output [7:0] mem_addr_out_137;            
  output [7:0] mem_addr_out_138;            
  output [7:0] mem_addr_out_139;            
  output [7:0] mem_addr_out_140;            
  output [7:0] mem_addr_out_141;            
  output [7:0] mem_addr_out_142;            
  output [7:0] mem_addr_out_143;            
  output [7:0] mem_addr_out_144;            
  output [7:0] mem_addr_out_145;            
  output [7:0] mem_addr_out_146;            
  output [7:0] mem_addr_out_147;            
  output [7:0] mem_addr_out_148;            
  output [7:0] mem_addr_out_149;            
  output [7:0] mem_addr_out_150;            
  output [7:0] mem_addr_out_151;            
  output [7:0] mem_addr_out_152;            
  output [7:0] mem_addr_out_153;            
  output [7:0] mem_addr_out_154;            
  output [7:0] mem_addr_out_155;            
  output [7:0] mem_addr_out_156;            
  output [7:0] mem_addr_out_157;            
  output [7:0] mem_addr_out_158;            
  output [7:0] mem_addr_out_159;            
  output [7:0] mem_addr_out_160;            
  output [7:0] mem_addr_out_161;            
  output [7:0] mem_addr_out_162;            
  output [7:0] mem_addr_out_163;            
  output [7:0] mem_addr_out_164;            
  output [7:0] mem_addr_out_165;            
  output [7:0] mem_addr_out_166;            
  output [7:0] mem_addr_out_167;            
  output [7:0] mem_addr_out_168;            
  output [7:0] mem_addr_out_169;            
  output [7:0] mem_addr_out_170;            
  output [7:0] mem_addr_out_171;            
  output [7:0] mem_addr_out_172;            
  output [7:0] mem_addr_out_173;            
  output [7:0] mem_addr_out_174;            
  output [7:0] mem_addr_out_175;            
  output [7:0] mem_addr_out_176;            
  output [7:0] mem_addr_out_177;            
  output [7:0] mem_addr_out_178;            
  output [7:0] mem_addr_out_179;            
  output [7:0] mem_addr_out_180;            
  output [7:0] mem_addr_out_181;            
  output [7:0] mem_addr_out_182;            
  output [7:0] mem_addr_out_183;            
  output [7:0] mem_addr_out_184;            
  output [7:0] mem_addr_out_185;            
  output [7:0] mem_addr_out_186;            
  output [7:0] mem_addr_out_187;            
  output [7:0] mem_addr_out_188;            
  output [7:0] mem_addr_out_189;            
  output [7:0] mem_addr_out_190;            
  output [7:0] mem_addr_out_191;            
  output [7:0] mem_addr_out_192;            
  output [7:0] mem_addr_out_193;            
  output [7:0] mem_addr_out_194;            
  output [7:0] mem_addr_out_195;            
  output [7:0] mem_addr_out_196;            
  output [7:0] mem_addr_out_197;            
  output [7:0] mem_addr_out_198;            
  output [7:0] mem_addr_out_199;            
  output [7:0] mem_addr_out_200;            
  output [7:0] mem_addr_out_201;            
  output [7:0] mem_addr_out_202;            
  output [7:0] mem_addr_out_203;            
  output [7:0] mem_addr_out_204;            
  output [7:0] mem_addr_out_205;            
  output [7:0] mem_addr_out_206;            
  output [7:0] mem_addr_out_207;            
  output [7:0] mem_addr_out_208;            
  output [7:0] mem_addr_out_209;            
  output [7:0] mem_addr_out_210;            
  output [7:0] mem_addr_out_211;            
  output [7:0] mem_addr_out_212;            
  output [7:0] mem_addr_out_213;            
  output [7:0] mem_addr_out_214;            
  output [7:0] mem_addr_out_215;            
  output [7:0] mem_addr_out_216;            
  output [7:0] mem_addr_out_217;            
  output [7:0] mem_addr_out_218;            
  output [7:0] mem_addr_out_219;            
  output [7:0] mem_addr_out_220;            
  output [7:0] mem_addr_out_221;            
  output [7:0] mem_addr_out_222;            
  output [7:0] mem_addr_out_223;            
  output [7:0] mem_addr_out_224;            
  output [7:0] mem_addr_out_225;            
  output [7:0] mem_addr_out_226;            
  output [7:0] mem_addr_out_227;            
  output [7:0] mem_addr_out_228;            
  output [7:0] mem_addr_out_229;            
  output [7:0] mem_addr_out_230;            
  output [7:0] mem_addr_out_231;            
  output [7:0] mem_addr_out_232;            
  output [7:0] mem_addr_out_233;            
  output [7:0] mem_addr_out_234;            
  output [7:0] mem_addr_out_235;            
  output [7:0] mem_addr_out_236;            
  output [7:0] mem_addr_out_237;            
  output [7:0] mem_addr_out_238;            
  output [7:0] mem_addr_out_239;            
  output [7:0] mem_addr_out_240;            
  output [7:0] mem_addr_out_241;            
  output [7:0] mem_addr_out_242;            
  output [7:0] mem_addr_out_243;            
  output [7:0] mem_addr_out_244;            
  output [7:0] mem_addr_out_245;            
  output [7:0] mem_addr_out_246;            
  output [7:0] mem_addr_out_247;            
  output [7:0] mem_addr_out_248;            
  output [7:0] mem_addr_out_249;            
  output [7:0] mem_addr_out_250;            
  output [7:0] mem_addr_out_251;            
  output [7:0] mem_addr_out_252;            
  output [7:0] mem_addr_out_253;            
  output [7:0] mem_addr_out_254;            
  output [7:0] mem_addr_out_255;            
  output wen_out;
  output reg out_start;
  
  reg [1:0] state;        
  reg flag;        

  wire [7:0] mem_addr_out_tmp_0;   
  wire [7:0] mem_addr_out_tmp_1;   
  wire [7:0] mem_addr_out_tmp_2;   
  wire [7:0] mem_addr_out_tmp_3;   
  wire [7:0] mem_addr_out_tmp_4;   
  wire [7:0] mem_addr_out_tmp_5;   
  wire [7:0] mem_addr_out_tmp_6;   
  wire [7:0] mem_addr_out_tmp_7;   
  wire [7:0] mem_addr_out_tmp_8;   
  wire [7:0] mem_addr_out_tmp_9;   
  wire [7:0] mem_addr_out_tmp_10;   
  wire [7:0] mem_addr_out_tmp_11;   
  wire [7:0] mem_addr_out_tmp_12;   
  wire [7:0] mem_addr_out_tmp_13;   
  wire [7:0] mem_addr_out_tmp_14;   
  wire [7:0] mem_addr_out_tmp_15;   
  wire [7:0] mem_addr_out_tmp_16;   
  wire [7:0] mem_addr_out_tmp_17;   
  wire [7:0] mem_addr_out_tmp_18;   
  wire [7:0] mem_addr_out_tmp_19;   
  wire [7:0] mem_addr_out_tmp_20;   
  wire [7:0] mem_addr_out_tmp_21;   
  wire [7:0] mem_addr_out_tmp_22;   
  wire [7:0] mem_addr_out_tmp_23;   
  wire [7:0] mem_addr_out_tmp_24;   
  wire [7:0] mem_addr_out_tmp_25;   
  wire [7:0] mem_addr_out_tmp_26;   
  wire [7:0] mem_addr_out_tmp_27;   
  wire [7:0] mem_addr_out_tmp_28;   
  wire [7:0] mem_addr_out_tmp_29;   
  wire [7:0] mem_addr_out_tmp_30;   
  wire [7:0] mem_addr_out_tmp_31;   
  wire [7:0] mem_addr_out_tmp_32;   
  wire [7:0] mem_addr_out_tmp_33;   
  wire [7:0] mem_addr_out_tmp_34;   
  wire [7:0] mem_addr_out_tmp_35;   
  wire [7:0] mem_addr_out_tmp_36;   
  wire [7:0] mem_addr_out_tmp_37;   
  wire [7:0] mem_addr_out_tmp_38;   
  wire [7:0] mem_addr_out_tmp_39;   
  wire [7:0] mem_addr_out_tmp_40;   
  wire [7:0] mem_addr_out_tmp_41;   
  wire [7:0] mem_addr_out_tmp_42;   
  wire [7:0] mem_addr_out_tmp_43;   
  wire [7:0] mem_addr_out_tmp_44;   
  wire [7:0] mem_addr_out_tmp_45;   
  wire [7:0] mem_addr_out_tmp_46;   
  wire [7:0] mem_addr_out_tmp_47;   
  wire [7:0] mem_addr_out_tmp_48;   
  wire [7:0] mem_addr_out_tmp_49;   
  wire [7:0] mem_addr_out_tmp_50;   
  wire [7:0] mem_addr_out_tmp_51;   
  wire [7:0] mem_addr_out_tmp_52;   
  wire [7:0] mem_addr_out_tmp_53;   
  wire [7:0] mem_addr_out_tmp_54;   
  wire [7:0] mem_addr_out_tmp_55;   
  wire [7:0] mem_addr_out_tmp_56;   
  wire [7:0] mem_addr_out_tmp_57;   
  wire [7:0] mem_addr_out_tmp_58;   
  wire [7:0] mem_addr_out_tmp_59;   
  wire [7:0] mem_addr_out_tmp_60;   
  wire [7:0] mem_addr_out_tmp_61;   
  wire [7:0] mem_addr_out_tmp_62;   
  wire [7:0] mem_addr_out_tmp_63;   
  wire [7:0] mem_addr_out_tmp_64;   
  wire [7:0] mem_addr_out_tmp_65;   
  wire [7:0] mem_addr_out_tmp_66;   
  wire [7:0] mem_addr_out_tmp_67;   
  wire [7:0] mem_addr_out_tmp_68;   
  wire [7:0] mem_addr_out_tmp_69;   
  wire [7:0] mem_addr_out_tmp_70;   
  wire [7:0] mem_addr_out_tmp_71;   
  wire [7:0] mem_addr_out_tmp_72;   
  wire [7:0] mem_addr_out_tmp_73;   
  wire [7:0] mem_addr_out_tmp_74;   
  wire [7:0] mem_addr_out_tmp_75;   
  wire [7:0] mem_addr_out_tmp_76;   
  wire [7:0] mem_addr_out_tmp_77;   
  wire [7:0] mem_addr_out_tmp_78;   
  wire [7:0] mem_addr_out_tmp_79;   
  wire [7:0] mem_addr_out_tmp_80;   
  wire [7:0] mem_addr_out_tmp_81;   
  wire [7:0] mem_addr_out_tmp_82;   
  wire [7:0] mem_addr_out_tmp_83;   
  wire [7:0] mem_addr_out_tmp_84;   
  wire [7:0] mem_addr_out_tmp_85;   
  wire [7:0] mem_addr_out_tmp_86;   
  wire [7:0] mem_addr_out_tmp_87;   
  wire [7:0] mem_addr_out_tmp_88;   
  wire [7:0] mem_addr_out_tmp_89;   
  wire [7:0] mem_addr_out_tmp_90;   
  wire [7:0] mem_addr_out_tmp_91;   
  wire [7:0] mem_addr_out_tmp_92;   
  wire [7:0] mem_addr_out_tmp_93;   
  wire [7:0] mem_addr_out_tmp_94;   
  wire [7:0] mem_addr_out_tmp_95;   
  wire [7:0] mem_addr_out_tmp_96;   
  wire [7:0] mem_addr_out_tmp_97;   
  wire [7:0] mem_addr_out_tmp_98;   
  wire [7:0] mem_addr_out_tmp_99;   
  wire [7:0] mem_addr_out_tmp_100;   
  wire [7:0] mem_addr_out_tmp_101;   
  wire [7:0] mem_addr_out_tmp_102;   
  wire [7:0] mem_addr_out_tmp_103;   
  wire [7:0] mem_addr_out_tmp_104;   
  wire [7:0] mem_addr_out_tmp_105;   
  wire [7:0] mem_addr_out_tmp_106;   
  wire [7:0] mem_addr_out_tmp_107;   
  wire [7:0] mem_addr_out_tmp_108;   
  wire [7:0] mem_addr_out_tmp_109;   
  wire [7:0] mem_addr_out_tmp_110;   
  wire [7:0] mem_addr_out_tmp_111;   
  wire [7:0] mem_addr_out_tmp_112;   
  wire [7:0] mem_addr_out_tmp_113;   
  wire [7:0] mem_addr_out_tmp_114;   
  wire [7:0] mem_addr_out_tmp_115;   
  wire [7:0] mem_addr_out_tmp_116;   
  wire [7:0] mem_addr_out_tmp_117;   
  wire [7:0] mem_addr_out_tmp_118;   
  wire [7:0] mem_addr_out_tmp_119;   
  wire [7:0] mem_addr_out_tmp_120;   
  wire [7:0] mem_addr_out_tmp_121;   
  wire [7:0] mem_addr_out_tmp_122;   
  wire [7:0] mem_addr_out_tmp_123;   
  wire [7:0] mem_addr_out_tmp_124;   
  wire [7:0] mem_addr_out_tmp_125;   
  wire [7:0] mem_addr_out_tmp_126;   
  wire [7:0] mem_addr_out_tmp_127;   
  wire [7:0] mem_addr_out_tmp_128;   
  wire [7:0] mem_addr_out_tmp_129;   
  wire [7:0] mem_addr_out_tmp_130;   
  wire [7:0] mem_addr_out_tmp_131;   
  wire [7:0] mem_addr_out_tmp_132;   
  wire [7:0] mem_addr_out_tmp_133;   
  wire [7:0] mem_addr_out_tmp_134;   
  wire [7:0] mem_addr_out_tmp_135;   
  wire [7:0] mem_addr_out_tmp_136;   
  wire [7:0] mem_addr_out_tmp_137;   
  wire [7:0] mem_addr_out_tmp_138;   
  wire [7:0] mem_addr_out_tmp_139;   
  wire [7:0] mem_addr_out_tmp_140;   
  wire [7:0] mem_addr_out_tmp_141;   
  wire [7:0] mem_addr_out_tmp_142;   
  wire [7:0] mem_addr_out_tmp_143;   
  wire [7:0] mem_addr_out_tmp_144;   
  wire [7:0] mem_addr_out_tmp_145;   
  wire [7:0] mem_addr_out_tmp_146;   
  wire [7:0] mem_addr_out_tmp_147;   
  wire [7:0] mem_addr_out_tmp_148;   
  wire [7:0] mem_addr_out_tmp_149;   
  wire [7:0] mem_addr_out_tmp_150;   
  wire [7:0] mem_addr_out_tmp_151;   
  wire [7:0] mem_addr_out_tmp_152;   
  wire [7:0] mem_addr_out_tmp_153;   
  wire [7:0] mem_addr_out_tmp_154;   
  wire [7:0] mem_addr_out_tmp_155;   
  wire [7:0] mem_addr_out_tmp_156;   
  wire [7:0] mem_addr_out_tmp_157;   
  wire [7:0] mem_addr_out_tmp_158;   
  wire [7:0] mem_addr_out_tmp_159;   
  wire [7:0] mem_addr_out_tmp_160;   
  wire [7:0] mem_addr_out_tmp_161;   
  wire [7:0] mem_addr_out_tmp_162;   
  wire [7:0] mem_addr_out_tmp_163;   
  wire [7:0] mem_addr_out_tmp_164;   
  wire [7:0] mem_addr_out_tmp_165;   
  wire [7:0] mem_addr_out_tmp_166;   
  wire [7:0] mem_addr_out_tmp_167;   
  wire [7:0] mem_addr_out_tmp_168;   
  wire [7:0] mem_addr_out_tmp_169;   
  wire [7:0] mem_addr_out_tmp_170;   
  wire [7:0] mem_addr_out_tmp_171;   
  wire [7:0] mem_addr_out_tmp_172;   
  wire [7:0] mem_addr_out_tmp_173;   
  wire [7:0] mem_addr_out_tmp_174;   
  wire [7:0] mem_addr_out_tmp_175;   
  wire [7:0] mem_addr_out_tmp_176;   
  wire [7:0] mem_addr_out_tmp_177;   
  wire [7:0] mem_addr_out_tmp_178;   
  wire [7:0] mem_addr_out_tmp_179;   
  wire [7:0] mem_addr_out_tmp_180;   
  wire [7:0] mem_addr_out_tmp_181;   
  wire [7:0] mem_addr_out_tmp_182;   
  wire [7:0] mem_addr_out_tmp_183;   
  wire [7:0] mem_addr_out_tmp_184;   
  wire [7:0] mem_addr_out_tmp_185;   
  wire [7:0] mem_addr_out_tmp_186;   
  wire [7:0] mem_addr_out_tmp_187;   
  wire [7:0] mem_addr_out_tmp_188;   
  wire [7:0] mem_addr_out_tmp_189;   
  wire [7:0] mem_addr_out_tmp_190;   
  wire [7:0] mem_addr_out_tmp_191;   
  wire [7:0] mem_addr_out_tmp_192;   
  wire [7:0] mem_addr_out_tmp_193;   
  wire [7:0] mem_addr_out_tmp_194;   
  wire [7:0] mem_addr_out_tmp_195;   
  wire [7:0] mem_addr_out_tmp_196;   
  wire [7:0] mem_addr_out_tmp_197;   
  wire [7:0] mem_addr_out_tmp_198;   
  wire [7:0] mem_addr_out_tmp_199;   
  wire [7:0] mem_addr_out_tmp_200;   
  wire [7:0] mem_addr_out_tmp_201;   
  wire [7:0] mem_addr_out_tmp_202;   
  wire [7:0] mem_addr_out_tmp_203;   
  wire [7:0] mem_addr_out_tmp_204;   
  wire [7:0] mem_addr_out_tmp_205;   
  wire [7:0] mem_addr_out_tmp_206;   
  wire [7:0] mem_addr_out_tmp_207;   
  wire [7:0] mem_addr_out_tmp_208;   
  wire [7:0] mem_addr_out_tmp_209;   
  wire [7:0] mem_addr_out_tmp_210;   
  wire [7:0] mem_addr_out_tmp_211;   
  wire [7:0] mem_addr_out_tmp_212;   
  wire [7:0] mem_addr_out_tmp_213;   
  wire [7:0] mem_addr_out_tmp_214;   
  wire [7:0] mem_addr_out_tmp_215;   
  wire [7:0] mem_addr_out_tmp_216;   
  wire [7:0] mem_addr_out_tmp_217;   
  wire [7:0] mem_addr_out_tmp_218;   
  wire [7:0] mem_addr_out_tmp_219;   
  wire [7:0] mem_addr_out_tmp_220;   
  wire [7:0] mem_addr_out_tmp_221;   
  wire [7:0] mem_addr_out_tmp_222;   
  wire [7:0] mem_addr_out_tmp_223;   
  wire [7:0] mem_addr_out_tmp_224;   
  wire [7:0] mem_addr_out_tmp_225;   
  wire [7:0] mem_addr_out_tmp_226;   
  wire [7:0] mem_addr_out_tmp_227;   
  wire [7:0] mem_addr_out_tmp_228;   
  wire [7:0] mem_addr_out_tmp_229;   
  wire [7:0] mem_addr_out_tmp_230;   
  wire [7:0] mem_addr_out_tmp_231;   
  wire [7:0] mem_addr_out_tmp_232;   
  wire [7:0] mem_addr_out_tmp_233;   
  wire [7:0] mem_addr_out_tmp_234;   
  wire [7:0] mem_addr_out_tmp_235;   
  wire [7:0] mem_addr_out_tmp_236;   
  wire [7:0] mem_addr_out_tmp_237;   
  wire [7:0] mem_addr_out_tmp_238;   
  wire [7:0] mem_addr_out_tmp_239;   
  wire [7:0] mem_addr_out_tmp_240;   
  wire [7:0] mem_addr_out_tmp_241;   
  wire [7:0] mem_addr_out_tmp_242;   
  wire [7:0] mem_addr_out_tmp_243;   
  wire [7:0] mem_addr_out_tmp_244;   
  wire [7:0] mem_addr_out_tmp_245;   
  wire [7:0] mem_addr_out_tmp_246;   
  wire [7:0] mem_addr_out_tmp_247;   
  wire [7:0] mem_addr_out_tmp_248;   
  wire [7:0] mem_addr_out_tmp_249;   
  wire [7:0] mem_addr_out_tmp_250;   
  wire [7:0] mem_addr_out_tmp_251;   
  wire [7:0] mem_addr_out_tmp_252;   
  wire [7:0] mem_addr_out_tmp_253;   
  wire [7:0] mem_addr_out_tmp_254;   
  wire [7:0] mem_addr_out_tmp_255;   
  wire [7:0] mem_addr_out_w;        
  wire [7:0] mem_addr_out_w_h;        
  
  mem_addr_gen_dp256_mem0_per0 top_mem_addr_gen_inst (.clk(clk),.rst(rst),.addr_out(mem_addr_out_w), .counter_in(counter_in)); 

  assign mem_addr_out_w_h = mem_addr_out_w[7:0];        
  assign mem_addr_out_tmp_0 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_1 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_2 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_3 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_4 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_5 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_6 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_7 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_8 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_9 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_10 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_11 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_12 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_13 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_14 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_15 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_16 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_17 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_18 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_19 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_20 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_21 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_22 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_23 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_24 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_25 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_26 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_27 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_28 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_29 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_30 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_31 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_32 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_33 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_34 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_35 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_36 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_37 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_38 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_39 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_40 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_41 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_42 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_43 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_44 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_45 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_46 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_47 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_48 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_49 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_50 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_51 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_52 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_53 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_54 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_55 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_56 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_57 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_58 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_59 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_60 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_61 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_62 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_63 = {mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_64 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_65 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_66 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_67 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_68 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_69 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_70 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_71 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_72 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_73 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_74 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_75 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_76 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_77 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_78 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_79 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_80 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_81 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_82 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_83 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_84 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_85 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_86 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_87 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_88 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_89 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_90 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_91 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_92 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_93 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_94 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_95 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_96 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_97 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_98 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_99 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_100 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_101 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_102 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_103 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_104 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_105 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_106 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_107 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_108 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_109 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_110 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_111 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_112 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_113 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_114 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_115 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_116 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_117 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_118 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_119 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_120 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_121 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_122 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_123 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_124 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_125 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_126 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_127 = {mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_128 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_129 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_130 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_131 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_132 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_133 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_134 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_135 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_136 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_137 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_138 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_139 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_140 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_141 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_142 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_143 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_144 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_145 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_146 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_147 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_148 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_149 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_150 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_151 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_152 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_153 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_154 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_155 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_156 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_157 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_158 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_159 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_160 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_161 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_162 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_163 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_164 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_165 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_166 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_167 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_168 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_169 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_170 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_171 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_172 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_173 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_174 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_175 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_176 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_177 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_178 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_179 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_180 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_181 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_182 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_183 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_184 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_185 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_186 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_187 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_188 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_189 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_190 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_191 = {~mem_addr_out_w_h[7],mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_192 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_193 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_194 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_195 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_196 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_197 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_198 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_199 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_200 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_201 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_202 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_203 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_204 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_205 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_206 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_207 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_208 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_209 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_210 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_211 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_212 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_213 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_214 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_215 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_216 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_217 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_218 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_219 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_220 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_221 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_222 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_223 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_224 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_225 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_226 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_227 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_228 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_229 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_230 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_231 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_232 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_233 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_234 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_235 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_236 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_237 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_238 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_239 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_240 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_241 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_242 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_243 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_244 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_245 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_246 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_247 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_248 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_249 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_250 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_251 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_252 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_253 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_254 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],mem_addr_out_w_h[0]}; 
  assign mem_addr_out_tmp_255 = {~mem_addr_out_w_h[7],~mem_addr_out_w_h[6],~mem_addr_out_w_h[5],~mem_addr_out_w_h[4],~mem_addr_out_w_h[3],~mem_addr_out_w_h[2],~mem_addr_out_w_h[1],~mem_addr_out_w_h[0]}; 
  assign mem_addr_out_0 = ((flag == 1'b0) ? mem_addr_out_tmp_0 : counter_in); 
  assign mem_addr_out_1 = ((flag == 1'b0) ? mem_addr_out_tmp_1 : counter_in); 
  assign mem_addr_out_2 = ((flag == 1'b0) ? mem_addr_out_tmp_2 : counter_in); 
  assign mem_addr_out_3 = ((flag == 1'b0) ? mem_addr_out_tmp_3 : counter_in); 
  assign mem_addr_out_4 = ((flag == 1'b0) ? mem_addr_out_tmp_4 : counter_in); 
  assign mem_addr_out_5 = ((flag == 1'b0) ? mem_addr_out_tmp_5 : counter_in); 
  assign mem_addr_out_6 = ((flag == 1'b0) ? mem_addr_out_tmp_6 : counter_in); 
  assign mem_addr_out_7 = ((flag == 1'b0) ? mem_addr_out_tmp_7 : counter_in); 
  assign mem_addr_out_8 = ((flag == 1'b0) ? mem_addr_out_tmp_8 : counter_in); 
  assign mem_addr_out_9 = ((flag == 1'b0) ? mem_addr_out_tmp_9 : counter_in); 
  assign mem_addr_out_10 = ((flag == 1'b0) ? mem_addr_out_tmp_10 : counter_in); 
  assign mem_addr_out_11 = ((flag == 1'b0) ? mem_addr_out_tmp_11 : counter_in); 
  assign mem_addr_out_12 = ((flag == 1'b0) ? mem_addr_out_tmp_12 : counter_in); 
  assign mem_addr_out_13 = ((flag == 1'b0) ? mem_addr_out_tmp_13 : counter_in); 
  assign mem_addr_out_14 = ((flag == 1'b0) ? mem_addr_out_tmp_14 : counter_in); 
  assign mem_addr_out_15 = ((flag == 1'b0) ? mem_addr_out_tmp_15 : counter_in); 
  assign mem_addr_out_16 = ((flag == 1'b0) ? mem_addr_out_tmp_16 : counter_in); 
  assign mem_addr_out_17 = ((flag == 1'b0) ? mem_addr_out_tmp_17 : counter_in); 
  assign mem_addr_out_18 = ((flag == 1'b0) ? mem_addr_out_tmp_18 : counter_in); 
  assign mem_addr_out_19 = ((flag == 1'b0) ? mem_addr_out_tmp_19 : counter_in); 
  assign mem_addr_out_20 = ((flag == 1'b0) ? mem_addr_out_tmp_20 : counter_in); 
  assign mem_addr_out_21 = ((flag == 1'b0) ? mem_addr_out_tmp_21 : counter_in); 
  assign mem_addr_out_22 = ((flag == 1'b0) ? mem_addr_out_tmp_22 : counter_in); 
  assign mem_addr_out_23 = ((flag == 1'b0) ? mem_addr_out_tmp_23 : counter_in); 
  assign mem_addr_out_24 = ((flag == 1'b0) ? mem_addr_out_tmp_24 : counter_in); 
  assign mem_addr_out_25 = ((flag == 1'b0) ? mem_addr_out_tmp_25 : counter_in); 
  assign mem_addr_out_26 = ((flag == 1'b0) ? mem_addr_out_tmp_26 : counter_in); 
  assign mem_addr_out_27 = ((flag == 1'b0) ? mem_addr_out_tmp_27 : counter_in); 
  assign mem_addr_out_28 = ((flag == 1'b0) ? mem_addr_out_tmp_28 : counter_in); 
  assign mem_addr_out_29 = ((flag == 1'b0) ? mem_addr_out_tmp_29 : counter_in); 
  assign mem_addr_out_30 = ((flag == 1'b0) ? mem_addr_out_tmp_30 : counter_in); 
  assign mem_addr_out_31 = ((flag == 1'b0) ? mem_addr_out_tmp_31 : counter_in); 
  assign mem_addr_out_32 = ((flag == 1'b0) ? mem_addr_out_tmp_32 : counter_in); 
  assign mem_addr_out_33 = ((flag == 1'b0) ? mem_addr_out_tmp_33 : counter_in); 
  assign mem_addr_out_34 = ((flag == 1'b0) ? mem_addr_out_tmp_34 : counter_in); 
  assign mem_addr_out_35 = ((flag == 1'b0) ? mem_addr_out_tmp_35 : counter_in); 
  assign mem_addr_out_36 = ((flag == 1'b0) ? mem_addr_out_tmp_36 : counter_in); 
  assign mem_addr_out_37 = ((flag == 1'b0) ? mem_addr_out_tmp_37 : counter_in); 
  assign mem_addr_out_38 = ((flag == 1'b0) ? mem_addr_out_tmp_38 : counter_in); 
  assign mem_addr_out_39 = ((flag == 1'b0) ? mem_addr_out_tmp_39 : counter_in); 
  assign mem_addr_out_40 = ((flag == 1'b0) ? mem_addr_out_tmp_40 : counter_in); 
  assign mem_addr_out_41 = ((flag == 1'b0) ? mem_addr_out_tmp_41 : counter_in); 
  assign mem_addr_out_42 = ((flag == 1'b0) ? mem_addr_out_tmp_42 : counter_in); 
  assign mem_addr_out_43 = ((flag == 1'b0) ? mem_addr_out_tmp_43 : counter_in); 
  assign mem_addr_out_44 = ((flag == 1'b0) ? mem_addr_out_tmp_44 : counter_in); 
  assign mem_addr_out_45 = ((flag == 1'b0) ? mem_addr_out_tmp_45 : counter_in); 
  assign mem_addr_out_46 = ((flag == 1'b0) ? mem_addr_out_tmp_46 : counter_in); 
  assign mem_addr_out_47 = ((flag == 1'b0) ? mem_addr_out_tmp_47 : counter_in); 
  assign mem_addr_out_48 = ((flag == 1'b0) ? mem_addr_out_tmp_48 : counter_in); 
  assign mem_addr_out_49 = ((flag == 1'b0) ? mem_addr_out_tmp_49 : counter_in); 
  assign mem_addr_out_50 = ((flag == 1'b0) ? mem_addr_out_tmp_50 : counter_in); 
  assign mem_addr_out_51 = ((flag == 1'b0) ? mem_addr_out_tmp_51 : counter_in); 
  assign mem_addr_out_52 = ((flag == 1'b0) ? mem_addr_out_tmp_52 : counter_in); 
  assign mem_addr_out_53 = ((flag == 1'b0) ? mem_addr_out_tmp_53 : counter_in); 
  assign mem_addr_out_54 = ((flag == 1'b0) ? mem_addr_out_tmp_54 : counter_in); 
  assign mem_addr_out_55 = ((flag == 1'b0) ? mem_addr_out_tmp_55 : counter_in); 
  assign mem_addr_out_56 = ((flag == 1'b0) ? mem_addr_out_tmp_56 : counter_in); 
  assign mem_addr_out_57 = ((flag == 1'b0) ? mem_addr_out_tmp_57 : counter_in); 
  assign mem_addr_out_58 = ((flag == 1'b0) ? mem_addr_out_tmp_58 : counter_in); 
  assign mem_addr_out_59 = ((flag == 1'b0) ? mem_addr_out_tmp_59 : counter_in); 
  assign mem_addr_out_60 = ((flag == 1'b0) ? mem_addr_out_tmp_60 : counter_in); 
  assign mem_addr_out_61 = ((flag == 1'b0) ? mem_addr_out_tmp_61 : counter_in); 
  assign mem_addr_out_62 = ((flag == 1'b0) ? mem_addr_out_tmp_62 : counter_in); 
  assign mem_addr_out_63 = ((flag == 1'b0) ? mem_addr_out_tmp_63 : counter_in); 
  assign mem_addr_out_64 = ((flag == 1'b0) ? mem_addr_out_tmp_64 : counter_in); 
  assign mem_addr_out_65 = ((flag == 1'b0) ? mem_addr_out_tmp_65 : counter_in); 
  assign mem_addr_out_66 = ((flag == 1'b0) ? mem_addr_out_tmp_66 : counter_in); 
  assign mem_addr_out_67 = ((flag == 1'b0) ? mem_addr_out_tmp_67 : counter_in); 
  assign mem_addr_out_68 = ((flag == 1'b0) ? mem_addr_out_tmp_68 : counter_in); 
  assign mem_addr_out_69 = ((flag == 1'b0) ? mem_addr_out_tmp_69 : counter_in); 
  assign mem_addr_out_70 = ((flag == 1'b0) ? mem_addr_out_tmp_70 : counter_in); 
  assign mem_addr_out_71 = ((flag == 1'b0) ? mem_addr_out_tmp_71 : counter_in); 
  assign mem_addr_out_72 = ((flag == 1'b0) ? mem_addr_out_tmp_72 : counter_in); 
  assign mem_addr_out_73 = ((flag == 1'b0) ? mem_addr_out_tmp_73 : counter_in); 
  assign mem_addr_out_74 = ((flag == 1'b0) ? mem_addr_out_tmp_74 : counter_in); 
  assign mem_addr_out_75 = ((flag == 1'b0) ? mem_addr_out_tmp_75 : counter_in); 
  assign mem_addr_out_76 = ((flag == 1'b0) ? mem_addr_out_tmp_76 : counter_in); 
  assign mem_addr_out_77 = ((flag == 1'b0) ? mem_addr_out_tmp_77 : counter_in); 
  assign mem_addr_out_78 = ((flag == 1'b0) ? mem_addr_out_tmp_78 : counter_in); 
  assign mem_addr_out_79 = ((flag == 1'b0) ? mem_addr_out_tmp_79 : counter_in); 
  assign mem_addr_out_80 = ((flag == 1'b0) ? mem_addr_out_tmp_80 : counter_in); 
  assign mem_addr_out_81 = ((flag == 1'b0) ? mem_addr_out_tmp_81 : counter_in); 
  assign mem_addr_out_82 = ((flag == 1'b0) ? mem_addr_out_tmp_82 : counter_in); 
  assign mem_addr_out_83 = ((flag == 1'b0) ? mem_addr_out_tmp_83 : counter_in); 
  assign mem_addr_out_84 = ((flag == 1'b0) ? mem_addr_out_tmp_84 : counter_in); 
  assign mem_addr_out_85 = ((flag == 1'b0) ? mem_addr_out_tmp_85 : counter_in); 
  assign mem_addr_out_86 = ((flag == 1'b0) ? mem_addr_out_tmp_86 : counter_in); 
  assign mem_addr_out_87 = ((flag == 1'b0) ? mem_addr_out_tmp_87 : counter_in); 
  assign mem_addr_out_88 = ((flag == 1'b0) ? mem_addr_out_tmp_88 : counter_in); 
  assign mem_addr_out_89 = ((flag == 1'b0) ? mem_addr_out_tmp_89 : counter_in); 
  assign mem_addr_out_90 = ((flag == 1'b0) ? mem_addr_out_tmp_90 : counter_in); 
  assign mem_addr_out_91 = ((flag == 1'b0) ? mem_addr_out_tmp_91 : counter_in); 
  assign mem_addr_out_92 = ((flag == 1'b0) ? mem_addr_out_tmp_92 : counter_in); 
  assign mem_addr_out_93 = ((flag == 1'b0) ? mem_addr_out_tmp_93 : counter_in); 
  assign mem_addr_out_94 = ((flag == 1'b0) ? mem_addr_out_tmp_94 : counter_in); 
  assign mem_addr_out_95 = ((flag == 1'b0) ? mem_addr_out_tmp_95 : counter_in); 
  assign mem_addr_out_96 = ((flag == 1'b0) ? mem_addr_out_tmp_96 : counter_in); 
  assign mem_addr_out_97 = ((flag == 1'b0) ? mem_addr_out_tmp_97 : counter_in); 
  assign mem_addr_out_98 = ((flag == 1'b0) ? mem_addr_out_tmp_98 : counter_in); 
  assign mem_addr_out_99 = ((flag == 1'b0) ? mem_addr_out_tmp_99 : counter_in); 
  assign mem_addr_out_100 = ((flag == 1'b0) ? mem_addr_out_tmp_100 : counter_in); 
  assign mem_addr_out_101 = ((flag == 1'b0) ? mem_addr_out_tmp_101 : counter_in); 
  assign mem_addr_out_102 = ((flag == 1'b0) ? mem_addr_out_tmp_102 : counter_in); 
  assign mem_addr_out_103 = ((flag == 1'b0) ? mem_addr_out_tmp_103 : counter_in); 
  assign mem_addr_out_104 = ((flag == 1'b0) ? mem_addr_out_tmp_104 : counter_in); 
  assign mem_addr_out_105 = ((flag == 1'b0) ? mem_addr_out_tmp_105 : counter_in); 
  assign mem_addr_out_106 = ((flag == 1'b0) ? mem_addr_out_tmp_106 : counter_in); 
  assign mem_addr_out_107 = ((flag == 1'b0) ? mem_addr_out_tmp_107 : counter_in); 
  assign mem_addr_out_108 = ((flag == 1'b0) ? mem_addr_out_tmp_108 : counter_in); 
  assign mem_addr_out_109 = ((flag == 1'b0) ? mem_addr_out_tmp_109 : counter_in); 
  assign mem_addr_out_110 = ((flag == 1'b0) ? mem_addr_out_tmp_110 : counter_in); 
  assign mem_addr_out_111 = ((flag == 1'b0) ? mem_addr_out_tmp_111 : counter_in); 
  assign mem_addr_out_112 = ((flag == 1'b0) ? mem_addr_out_tmp_112 : counter_in); 
  assign mem_addr_out_113 = ((flag == 1'b0) ? mem_addr_out_tmp_113 : counter_in); 
  assign mem_addr_out_114 = ((flag == 1'b0) ? mem_addr_out_tmp_114 : counter_in); 
  assign mem_addr_out_115 = ((flag == 1'b0) ? mem_addr_out_tmp_115 : counter_in); 
  assign mem_addr_out_116 = ((flag == 1'b0) ? mem_addr_out_tmp_116 : counter_in); 
  assign mem_addr_out_117 = ((flag == 1'b0) ? mem_addr_out_tmp_117 : counter_in); 
  assign mem_addr_out_118 = ((flag == 1'b0) ? mem_addr_out_tmp_118 : counter_in); 
  assign mem_addr_out_119 = ((flag == 1'b0) ? mem_addr_out_tmp_119 : counter_in); 
  assign mem_addr_out_120 = ((flag == 1'b0) ? mem_addr_out_tmp_120 : counter_in); 
  assign mem_addr_out_121 = ((flag == 1'b0) ? mem_addr_out_tmp_121 : counter_in); 
  assign mem_addr_out_122 = ((flag == 1'b0) ? mem_addr_out_tmp_122 : counter_in); 
  assign mem_addr_out_123 = ((flag == 1'b0) ? mem_addr_out_tmp_123 : counter_in); 
  assign mem_addr_out_124 = ((flag == 1'b0) ? mem_addr_out_tmp_124 : counter_in); 
  assign mem_addr_out_125 = ((flag == 1'b0) ? mem_addr_out_tmp_125 : counter_in); 
  assign mem_addr_out_126 = ((flag == 1'b0) ? mem_addr_out_tmp_126 : counter_in); 
  assign mem_addr_out_127 = ((flag == 1'b0) ? mem_addr_out_tmp_127 : counter_in); 
  assign mem_addr_out_128 = ((flag == 1'b0) ? mem_addr_out_tmp_128 : counter_in); 
  assign mem_addr_out_129 = ((flag == 1'b0) ? mem_addr_out_tmp_129 : counter_in); 
  assign mem_addr_out_130 = ((flag == 1'b0) ? mem_addr_out_tmp_130 : counter_in); 
  assign mem_addr_out_131 = ((flag == 1'b0) ? mem_addr_out_tmp_131 : counter_in); 
  assign mem_addr_out_132 = ((flag == 1'b0) ? mem_addr_out_tmp_132 : counter_in); 
  assign mem_addr_out_133 = ((flag == 1'b0) ? mem_addr_out_tmp_133 : counter_in); 
  assign mem_addr_out_134 = ((flag == 1'b0) ? mem_addr_out_tmp_134 : counter_in); 
  assign mem_addr_out_135 = ((flag == 1'b0) ? mem_addr_out_tmp_135 : counter_in); 
  assign mem_addr_out_136 = ((flag == 1'b0) ? mem_addr_out_tmp_136 : counter_in); 
  assign mem_addr_out_137 = ((flag == 1'b0) ? mem_addr_out_tmp_137 : counter_in); 
  assign mem_addr_out_138 = ((flag == 1'b0) ? mem_addr_out_tmp_138 : counter_in); 
  assign mem_addr_out_139 = ((flag == 1'b0) ? mem_addr_out_tmp_139 : counter_in); 
  assign mem_addr_out_140 = ((flag == 1'b0) ? mem_addr_out_tmp_140 : counter_in); 
  assign mem_addr_out_141 = ((flag == 1'b0) ? mem_addr_out_tmp_141 : counter_in); 
  assign mem_addr_out_142 = ((flag == 1'b0) ? mem_addr_out_tmp_142 : counter_in); 
  assign mem_addr_out_143 = ((flag == 1'b0) ? mem_addr_out_tmp_143 : counter_in); 
  assign mem_addr_out_144 = ((flag == 1'b0) ? mem_addr_out_tmp_144 : counter_in); 
  assign mem_addr_out_145 = ((flag == 1'b0) ? mem_addr_out_tmp_145 : counter_in); 
  assign mem_addr_out_146 = ((flag == 1'b0) ? mem_addr_out_tmp_146 : counter_in); 
  assign mem_addr_out_147 = ((flag == 1'b0) ? mem_addr_out_tmp_147 : counter_in); 
  assign mem_addr_out_148 = ((flag == 1'b0) ? mem_addr_out_tmp_148 : counter_in); 
  assign mem_addr_out_149 = ((flag == 1'b0) ? mem_addr_out_tmp_149 : counter_in); 
  assign mem_addr_out_150 = ((flag == 1'b0) ? mem_addr_out_tmp_150 : counter_in); 
  assign mem_addr_out_151 = ((flag == 1'b0) ? mem_addr_out_tmp_151 : counter_in); 
  assign mem_addr_out_152 = ((flag == 1'b0) ? mem_addr_out_tmp_152 : counter_in); 
  assign mem_addr_out_153 = ((flag == 1'b0) ? mem_addr_out_tmp_153 : counter_in); 
  assign mem_addr_out_154 = ((flag == 1'b0) ? mem_addr_out_tmp_154 : counter_in); 
  assign mem_addr_out_155 = ((flag == 1'b0) ? mem_addr_out_tmp_155 : counter_in); 
  assign mem_addr_out_156 = ((flag == 1'b0) ? mem_addr_out_tmp_156 : counter_in); 
  assign mem_addr_out_157 = ((flag == 1'b0) ? mem_addr_out_tmp_157 : counter_in); 
  assign mem_addr_out_158 = ((flag == 1'b0) ? mem_addr_out_tmp_158 : counter_in); 
  assign mem_addr_out_159 = ((flag == 1'b0) ? mem_addr_out_tmp_159 : counter_in); 
  assign mem_addr_out_160 = ((flag == 1'b0) ? mem_addr_out_tmp_160 : counter_in); 
  assign mem_addr_out_161 = ((flag == 1'b0) ? mem_addr_out_tmp_161 : counter_in); 
  assign mem_addr_out_162 = ((flag == 1'b0) ? mem_addr_out_tmp_162 : counter_in); 
  assign mem_addr_out_163 = ((flag == 1'b0) ? mem_addr_out_tmp_163 : counter_in); 
  assign mem_addr_out_164 = ((flag == 1'b0) ? mem_addr_out_tmp_164 : counter_in); 
  assign mem_addr_out_165 = ((flag == 1'b0) ? mem_addr_out_tmp_165 : counter_in); 
  assign mem_addr_out_166 = ((flag == 1'b0) ? mem_addr_out_tmp_166 : counter_in); 
  assign mem_addr_out_167 = ((flag == 1'b0) ? mem_addr_out_tmp_167 : counter_in); 
  assign mem_addr_out_168 = ((flag == 1'b0) ? mem_addr_out_tmp_168 : counter_in); 
  assign mem_addr_out_169 = ((flag == 1'b0) ? mem_addr_out_tmp_169 : counter_in); 
  assign mem_addr_out_170 = ((flag == 1'b0) ? mem_addr_out_tmp_170 : counter_in); 
  assign mem_addr_out_171 = ((flag == 1'b0) ? mem_addr_out_tmp_171 : counter_in); 
  assign mem_addr_out_172 = ((flag == 1'b0) ? mem_addr_out_tmp_172 : counter_in); 
  assign mem_addr_out_173 = ((flag == 1'b0) ? mem_addr_out_tmp_173 : counter_in); 
  assign mem_addr_out_174 = ((flag == 1'b0) ? mem_addr_out_tmp_174 : counter_in); 
  assign mem_addr_out_175 = ((flag == 1'b0) ? mem_addr_out_tmp_175 : counter_in); 
  assign mem_addr_out_176 = ((flag == 1'b0) ? mem_addr_out_tmp_176 : counter_in); 
  assign mem_addr_out_177 = ((flag == 1'b0) ? mem_addr_out_tmp_177 : counter_in); 
  assign mem_addr_out_178 = ((flag == 1'b0) ? mem_addr_out_tmp_178 : counter_in); 
  assign mem_addr_out_179 = ((flag == 1'b0) ? mem_addr_out_tmp_179 : counter_in); 
  assign mem_addr_out_180 = ((flag == 1'b0) ? mem_addr_out_tmp_180 : counter_in); 
  assign mem_addr_out_181 = ((flag == 1'b0) ? mem_addr_out_tmp_181 : counter_in); 
  assign mem_addr_out_182 = ((flag == 1'b0) ? mem_addr_out_tmp_182 : counter_in); 
  assign mem_addr_out_183 = ((flag == 1'b0) ? mem_addr_out_tmp_183 : counter_in); 
  assign mem_addr_out_184 = ((flag == 1'b0) ? mem_addr_out_tmp_184 : counter_in); 
  assign mem_addr_out_185 = ((flag == 1'b0) ? mem_addr_out_tmp_185 : counter_in); 
  assign mem_addr_out_186 = ((flag == 1'b0) ? mem_addr_out_tmp_186 : counter_in); 
  assign mem_addr_out_187 = ((flag == 1'b0) ? mem_addr_out_tmp_187 : counter_in); 
  assign mem_addr_out_188 = ((flag == 1'b0) ? mem_addr_out_tmp_188 : counter_in); 
  assign mem_addr_out_189 = ((flag == 1'b0) ? mem_addr_out_tmp_189 : counter_in); 
  assign mem_addr_out_190 = ((flag == 1'b0) ? mem_addr_out_tmp_190 : counter_in); 
  assign mem_addr_out_191 = ((flag == 1'b0) ? mem_addr_out_tmp_191 : counter_in); 
  assign mem_addr_out_192 = ((flag == 1'b0) ? mem_addr_out_tmp_192 : counter_in); 
  assign mem_addr_out_193 = ((flag == 1'b0) ? mem_addr_out_tmp_193 : counter_in); 
  assign mem_addr_out_194 = ((flag == 1'b0) ? mem_addr_out_tmp_194 : counter_in); 
  assign mem_addr_out_195 = ((flag == 1'b0) ? mem_addr_out_tmp_195 : counter_in); 
  assign mem_addr_out_196 = ((flag == 1'b0) ? mem_addr_out_tmp_196 : counter_in); 
  assign mem_addr_out_197 = ((flag == 1'b0) ? mem_addr_out_tmp_197 : counter_in); 
  assign mem_addr_out_198 = ((flag == 1'b0) ? mem_addr_out_tmp_198 : counter_in); 
  assign mem_addr_out_199 = ((flag == 1'b0) ? mem_addr_out_tmp_199 : counter_in); 
  assign mem_addr_out_200 = ((flag == 1'b0) ? mem_addr_out_tmp_200 : counter_in); 
  assign mem_addr_out_201 = ((flag == 1'b0) ? mem_addr_out_tmp_201 : counter_in); 
  assign mem_addr_out_202 = ((flag == 1'b0) ? mem_addr_out_tmp_202 : counter_in); 
  assign mem_addr_out_203 = ((flag == 1'b0) ? mem_addr_out_tmp_203 : counter_in); 
  assign mem_addr_out_204 = ((flag == 1'b0) ? mem_addr_out_tmp_204 : counter_in); 
  assign mem_addr_out_205 = ((flag == 1'b0) ? mem_addr_out_tmp_205 : counter_in); 
  assign mem_addr_out_206 = ((flag == 1'b0) ? mem_addr_out_tmp_206 : counter_in); 
  assign mem_addr_out_207 = ((flag == 1'b0) ? mem_addr_out_tmp_207 : counter_in); 
  assign mem_addr_out_208 = ((flag == 1'b0) ? mem_addr_out_tmp_208 : counter_in); 
  assign mem_addr_out_209 = ((flag == 1'b0) ? mem_addr_out_tmp_209 : counter_in); 
  assign mem_addr_out_210 = ((flag == 1'b0) ? mem_addr_out_tmp_210 : counter_in); 
  assign mem_addr_out_211 = ((flag == 1'b0) ? mem_addr_out_tmp_211 : counter_in); 
  assign mem_addr_out_212 = ((flag == 1'b0) ? mem_addr_out_tmp_212 : counter_in); 
  assign mem_addr_out_213 = ((flag == 1'b0) ? mem_addr_out_tmp_213 : counter_in); 
  assign mem_addr_out_214 = ((flag == 1'b0) ? mem_addr_out_tmp_214 : counter_in); 
  assign mem_addr_out_215 = ((flag == 1'b0) ? mem_addr_out_tmp_215 : counter_in); 
  assign mem_addr_out_216 = ((flag == 1'b0) ? mem_addr_out_tmp_216 : counter_in); 
  assign mem_addr_out_217 = ((flag == 1'b0) ? mem_addr_out_tmp_217 : counter_in); 
  assign mem_addr_out_218 = ((flag == 1'b0) ? mem_addr_out_tmp_218 : counter_in); 
  assign mem_addr_out_219 = ((flag == 1'b0) ? mem_addr_out_tmp_219 : counter_in); 
  assign mem_addr_out_220 = ((flag == 1'b0) ? mem_addr_out_tmp_220 : counter_in); 
  assign mem_addr_out_221 = ((flag == 1'b0) ? mem_addr_out_tmp_221 : counter_in); 
  assign mem_addr_out_222 = ((flag == 1'b0) ? mem_addr_out_tmp_222 : counter_in); 
  assign mem_addr_out_223 = ((flag == 1'b0) ? mem_addr_out_tmp_223 : counter_in); 
  assign mem_addr_out_224 = ((flag == 1'b0) ? mem_addr_out_tmp_224 : counter_in); 
  assign mem_addr_out_225 = ((flag == 1'b0) ? mem_addr_out_tmp_225 : counter_in); 
  assign mem_addr_out_226 = ((flag == 1'b0) ? mem_addr_out_tmp_226 : counter_in); 
  assign mem_addr_out_227 = ((flag == 1'b0) ? mem_addr_out_tmp_227 : counter_in); 
  assign mem_addr_out_228 = ((flag == 1'b0) ? mem_addr_out_tmp_228 : counter_in); 
  assign mem_addr_out_229 = ((flag == 1'b0) ? mem_addr_out_tmp_229 : counter_in); 
  assign mem_addr_out_230 = ((flag == 1'b0) ? mem_addr_out_tmp_230 : counter_in); 
  assign mem_addr_out_231 = ((flag == 1'b0) ? mem_addr_out_tmp_231 : counter_in); 
  assign mem_addr_out_232 = ((flag == 1'b0) ? mem_addr_out_tmp_232 : counter_in); 
  assign mem_addr_out_233 = ((flag == 1'b0) ? mem_addr_out_tmp_233 : counter_in); 
  assign mem_addr_out_234 = ((flag == 1'b0) ? mem_addr_out_tmp_234 : counter_in); 
  assign mem_addr_out_235 = ((flag == 1'b0) ? mem_addr_out_tmp_235 : counter_in); 
  assign mem_addr_out_236 = ((flag == 1'b0) ? mem_addr_out_tmp_236 : counter_in); 
  assign mem_addr_out_237 = ((flag == 1'b0) ? mem_addr_out_tmp_237 : counter_in); 
  assign mem_addr_out_238 = ((flag == 1'b0) ? mem_addr_out_tmp_238 : counter_in); 
  assign mem_addr_out_239 = ((flag == 1'b0) ? mem_addr_out_tmp_239 : counter_in); 
  assign mem_addr_out_240 = ((flag == 1'b0) ? mem_addr_out_tmp_240 : counter_in); 
  assign mem_addr_out_241 = ((flag == 1'b0) ? mem_addr_out_tmp_241 : counter_in); 
  assign mem_addr_out_242 = ((flag == 1'b0) ? mem_addr_out_tmp_242 : counter_in); 
  assign mem_addr_out_243 = ((flag == 1'b0) ? mem_addr_out_tmp_243 : counter_in); 
  assign mem_addr_out_244 = ((flag == 1'b0) ? mem_addr_out_tmp_244 : counter_in); 
  assign mem_addr_out_245 = ((flag == 1'b0) ? mem_addr_out_tmp_245 : counter_in); 
  assign mem_addr_out_246 = ((flag == 1'b0) ? mem_addr_out_tmp_246 : counter_in); 
  assign mem_addr_out_247 = ((flag == 1'b0) ? mem_addr_out_tmp_247 : counter_in); 
  assign mem_addr_out_248 = ((flag == 1'b0) ? mem_addr_out_tmp_248 : counter_in); 
  assign mem_addr_out_249 = ((flag == 1'b0) ? mem_addr_out_tmp_249 : counter_in); 
  assign mem_addr_out_250 = ((flag == 1'b0) ? mem_addr_out_tmp_250 : counter_in); 
  assign mem_addr_out_251 = ((flag == 1'b0) ? mem_addr_out_tmp_251 : counter_in); 
  assign mem_addr_out_252 = ((flag == 1'b0) ? mem_addr_out_tmp_252 : counter_in); 
  assign mem_addr_out_253 = ((flag == 1'b0) ? mem_addr_out_tmp_253 : counter_in); 
  assign mem_addr_out_254 = ((flag == 1'b0) ? mem_addr_out_tmp_254 : counter_in); 
  assign mem_addr_out_255 = ((flag == 1'b0) ? mem_addr_out_tmp_255 : counter_in); 
  
  assign wen_out = state[0];        
  always@(posedge clk)             
  begin                            
    if(rst) begin                    
      out_start <= 1'b0; 
end
    else begin                        
      out_start <= (state == 2'b01) && (counter_in[7:0] == {8{1'b1}}); 
end                              
end                              

  always@(posedge clk)             
  begin                            
    if(rst) begin                    
      state <= 2'b0;            
      flag <= 1'b0;            
      end
    else begin                        
      case (state)              
        2'b00: begin              
          if (in_start)  begin              
            state <= 2'b01;              
            end
        end
        2'b01: begin              
          if (!in_start && counter_in == {8{1'b1}})  begin 
            state <= 2'b11;              
          end
          if (counter_in == {8{1'b1}})  begin 
            flag <= !flag;              
          end
        end
        2'b11: begin              
          if (counter_in == {8{1'b1}})  begin 
            state <= 2'b00;              
          end
        end
        default: state <= 2'b00;       
      endcase
    end
  end                              

endmodule                        


module mem_stage_dp256_r(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
clk,                             
counter_in,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;                   
  input [8-1:0] counter_in;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output reg [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255;
  output reg out_start; 
  
  wire [DATA_WIDTH-1:0] wire_in [255:0];              
  wire [DATA_WIDTH-1:0] wire_out [255:0];              
  
  wire wen_wire;              
  wire out_start_wire;              
  assign wire_in[0] = inData_0;    
  assign wire_in[1] = inData_1;    
  assign wire_in[2] = inData_2;    
  assign wire_in[3] = inData_3;    
  assign wire_in[4] = inData_4;    
  assign wire_in[5] = inData_5;    
  assign wire_in[6] = inData_6;    
  assign wire_in[7] = inData_7;    
  assign wire_in[8] = inData_8;    
  assign wire_in[9] = inData_9;    
  assign wire_in[10] = inData_10;    
  assign wire_in[11] = inData_11;    
  assign wire_in[12] = inData_12;    
  assign wire_in[13] = inData_13;    
  assign wire_in[14] = inData_14;    
  assign wire_in[15] = inData_15;    
  assign wire_in[16] = inData_16;    
  assign wire_in[17] = inData_17;    
  assign wire_in[18] = inData_18;    
  assign wire_in[19] = inData_19;    
  assign wire_in[20] = inData_20;    
  assign wire_in[21] = inData_21;    
  assign wire_in[22] = inData_22;    
  assign wire_in[23] = inData_23;    
  assign wire_in[24] = inData_24;    
  assign wire_in[25] = inData_25;    
  assign wire_in[26] = inData_26;    
  assign wire_in[27] = inData_27;    
  assign wire_in[28] = inData_28;    
  assign wire_in[29] = inData_29;    
  assign wire_in[30] = inData_30;    
  assign wire_in[31] = inData_31;    
  assign wire_in[32] = inData_32;    
  assign wire_in[33] = inData_33;    
  assign wire_in[34] = inData_34;    
  assign wire_in[35] = inData_35;    
  assign wire_in[36] = inData_36;    
  assign wire_in[37] = inData_37;    
  assign wire_in[38] = inData_38;    
  assign wire_in[39] = inData_39;    
  assign wire_in[40] = inData_40;    
  assign wire_in[41] = inData_41;    
  assign wire_in[42] = inData_42;    
  assign wire_in[43] = inData_43;    
  assign wire_in[44] = inData_44;    
  assign wire_in[45] = inData_45;    
  assign wire_in[46] = inData_46;    
  assign wire_in[47] = inData_47;    
  assign wire_in[48] = inData_48;    
  assign wire_in[49] = inData_49;    
  assign wire_in[50] = inData_50;    
  assign wire_in[51] = inData_51;    
  assign wire_in[52] = inData_52;    
  assign wire_in[53] = inData_53;    
  assign wire_in[54] = inData_54;    
  assign wire_in[55] = inData_55;    
  assign wire_in[56] = inData_56;    
  assign wire_in[57] = inData_57;    
  assign wire_in[58] = inData_58;    
  assign wire_in[59] = inData_59;    
  assign wire_in[60] = inData_60;    
  assign wire_in[61] = inData_61;    
  assign wire_in[62] = inData_62;    
  assign wire_in[63] = inData_63;    
  assign wire_in[64] = inData_64;    
  assign wire_in[65] = inData_65;    
  assign wire_in[66] = inData_66;    
  assign wire_in[67] = inData_67;    
  assign wire_in[68] = inData_68;    
  assign wire_in[69] = inData_69;    
  assign wire_in[70] = inData_70;    
  assign wire_in[71] = inData_71;    
  assign wire_in[72] = inData_72;    
  assign wire_in[73] = inData_73;    
  assign wire_in[74] = inData_74;    
  assign wire_in[75] = inData_75;    
  assign wire_in[76] = inData_76;    
  assign wire_in[77] = inData_77;    
  assign wire_in[78] = inData_78;    
  assign wire_in[79] = inData_79;    
  assign wire_in[80] = inData_80;    
  assign wire_in[81] = inData_81;    
  assign wire_in[82] = inData_82;    
  assign wire_in[83] = inData_83;    
  assign wire_in[84] = inData_84;    
  assign wire_in[85] = inData_85;    
  assign wire_in[86] = inData_86;    
  assign wire_in[87] = inData_87;    
  assign wire_in[88] = inData_88;    
  assign wire_in[89] = inData_89;    
  assign wire_in[90] = inData_90;    
  assign wire_in[91] = inData_91;    
  assign wire_in[92] = inData_92;    
  assign wire_in[93] = inData_93;    
  assign wire_in[94] = inData_94;    
  assign wire_in[95] = inData_95;    
  assign wire_in[96] = inData_96;    
  assign wire_in[97] = inData_97;    
  assign wire_in[98] = inData_98;    
  assign wire_in[99] = inData_99;    
  assign wire_in[100] = inData_100;    
  assign wire_in[101] = inData_101;    
  assign wire_in[102] = inData_102;    
  assign wire_in[103] = inData_103;    
  assign wire_in[104] = inData_104;    
  assign wire_in[105] = inData_105;    
  assign wire_in[106] = inData_106;    
  assign wire_in[107] = inData_107;    
  assign wire_in[108] = inData_108;    
  assign wire_in[109] = inData_109;    
  assign wire_in[110] = inData_110;    
  assign wire_in[111] = inData_111;    
  assign wire_in[112] = inData_112;    
  assign wire_in[113] = inData_113;    
  assign wire_in[114] = inData_114;    
  assign wire_in[115] = inData_115;    
  assign wire_in[116] = inData_116;    
  assign wire_in[117] = inData_117;    
  assign wire_in[118] = inData_118;    
  assign wire_in[119] = inData_119;    
  assign wire_in[120] = inData_120;    
  assign wire_in[121] = inData_121;    
  assign wire_in[122] = inData_122;    
  assign wire_in[123] = inData_123;    
  assign wire_in[124] = inData_124;    
  assign wire_in[125] = inData_125;    
  assign wire_in[126] = inData_126;    
  assign wire_in[127] = inData_127;    
  assign wire_in[128] = inData_128;    
  assign wire_in[129] = inData_129;    
  assign wire_in[130] = inData_130;    
  assign wire_in[131] = inData_131;    
  assign wire_in[132] = inData_132;    
  assign wire_in[133] = inData_133;    
  assign wire_in[134] = inData_134;    
  assign wire_in[135] = inData_135;    
  assign wire_in[136] = inData_136;    
  assign wire_in[137] = inData_137;    
  assign wire_in[138] = inData_138;    
  assign wire_in[139] = inData_139;    
  assign wire_in[140] = inData_140;    
  assign wire_in[141] = inData_141;    
  assign wire_in[142] = inData_142;    
  assign wire_in[143] = inData_143;    
  assign wire_in[144] = inData_144;    
  assign wire_in[145] = inData_145;    
  assign wire_in[146] = inData_146;    
  assign wire_in[147] = inData_147;    
  assign wire_in[148] = inData_148;    
  assign wire_in[149] = inData_149;    
  assign wire_in[150] = inData_150;    
  assign wire_in[151] = inData_151;    
  assign wire_in[152] = inData_152;    
  assign wire_in[153] = inData_153;    
  assign wire_in[154] = inData_154;    
  assign wire_in[155] = inData_155;    
  assign wire_in[156] = inData_156;    
  assign wire_in[157] = inData_157;    
  assign wire_in[158] = inData_158;    
  assign wire_in[159] = inData_159;    
  assign wire_in[160] = inData_160;    
  assign wire_in[161] = inData_161;    
  assign wire_in[162] = inData_162;    
  assign wire_in[163] = inData_163;    
  assign wire_in[164] = inData_164;    
  assign wire_in[165] = inData_165;    
  assign wire_in[166] = inData_166;    
  assign wire_in[167] = inData_167;    
  assign wire_in[168] = inData_168;    
  assign wire_in[169] = inData_169;    
  assign wire_in[170] = inData_170;    
  assign wire_in[171] = inData_171;    
  assign wire_in[172] = inData_172;    
  assign wire_in[173] = inData_173;    
  assign wire_in[174] = inData_174;    
  assign wire_in[175] = inData_175;    
  assign wire_in[176] = inData_176;    
  assign wire_in[177] = inData_177;    
  assign wire_in[178] = inData_178;    
  assign wire_in[179] = inData_179;    
  assign wire_in[180] = inData_180;    
  assign wire_in[181] = inData_181;    
  assign wire_in[182] = inData_182;    
  assign wire_in[183] = inData_183;    
  assign wire_in[184] = inData_184;    
  assign wire_in[185] = inData_185;    
  assign wire_in[186] = inData_186;    
  assign wire_in[187] = inData_187;    
  assign wire_in[188] = inData_188;    
  assign wire_in[189] = inData_189;    
  assign wire_in[190] = inData_190;    
  assign wire_in[191] = inData_191;    
  assign wire_in[192] = inData_192;    
  assign wire_in[193] = inData_193;    
  assign wire_in[194] = inData_194;    
  assign wire_in[195] = inData_195;    
  assign wire_in[196] = inData_196;    
  assign wire_in[197] = inData_197;    
  assign wire_in[198] = inData_198;    
  assign wire_in[199] = inData_199;    
  assign wire_in[200] = inData_200;    
  assign wire_in[201] = inData_201;    
  assign wire_in[202] = inData_202;    
  assign wire_in[203] = inData_203;    
  assign wire_in[204] = inData_204;    
  assign wire_in[205] = inData_205;    
  assign wire_in[206] = inData_206;    
  assign wire_in[207] = inData_207;    
  assign wire_in[208] = inData_208;    
  assign wire_in[209] = inData_209;    
  assign wire_in[210] = inData_210;    
  assign wire_in[211] = inData_211;    
  assign wire_in[212] = inData_212;    
  assign wire_in[213] = inData_213;    
  assign wire_in[214] = inData_214;    
  assign wire_in[215] = inData_215;    
  assign wire_in[216] = inData_216;    
  assign wire_in[217] = inData_217;    
  assign wire_in[218] = inData_218;    
  assign wire_in[219] = inData_219;    
  assign wire_in[220] = inData_220;    
  assign wire_in[221] = inData_221;    
  assign wire_in[222] = inData_222;    
  assign wire_in[223] = inData_223;    
  assign wire_in[224] = inData_224;    
  assign wire_in[225] = inData_225;    
  assign wire_in[226] = inData_226;    
  assign wire_in[227] = inData_227;    
  assign wire_in[228] = inData_228;    
  assign wire_in[229] = inData_229;    
  assign wire_in[230] = inData_230;    
  assign wire_in[231] = inData_231;    
  assign wire_in[232] = inData_232;    
  assign wire_in[233] = inData_233;    
  assign wire_in[234] = inData_234;    
  assign wire_in[235] = inData_235;    
  assign wire_in[236] = inData_236;    
  assign wire_in[237] = inData_237;    
  assign wire_in[238] = inData_238;    
  assign wire_in[239] = inData_239;    
  assign wire_in[240] = inData_240;    
  assign wire_in[241] = inData_241;    
  assign wire_in[242] = inData_242;    
  assign wire_in[243] = inData_243;    
  assign wire_in[244] = inData_244;    
  assign wire_in[245] = inData_245;    
  assign wire_in[246] = inData_246;    
  assign wire_in[247] = inData_247;    
  assign wire_in[248] = inData_248;    
  assign wire_in[249] = inData_249;    
  assign wire_in[250] = inData_250;    
  assign wire_in[251] = inData_251;    
  assign wire_in[252] = inData_252;    
  assign wire_in[253] = inData_253;    
  assign wire_in[254] = inData_254;    
  assign wire_in[255] = inData_255;    
  
  wire [7:0] addr_w_wire_0;        

  wire [7:0] addr_w_wire_1;        

  wire [7:0] addr_w_wire_2;        

  wire [7:0] addr_w_wire_3;        

  wire [7:0] addr_w_wire_4;        

  wire [7:0] addr_w_wire_5;        

  wire [7:0] addr_w_wire_6;        

  wire [7:0] addr_w_wire_7;        

  wire [7:0] addr_w_wire_8;        

  wire [7:0] addr_w_wire_9;        

  wire [7:0] addr_w_wire_10;        

  wire [7:0] addr_w_wire_11;        

  wire [7:0] addr_w_wire_12;        

  wire [7:0] addr_w_wire_13;        

  wire [7:0] addr_w_wire_14;        

  wire [7:0] addr_w_wire_15;        

  wire [7:0] addr_w_wire_16;        

  wire [7:0] addr_w_wire_17;        

  wire [7:0] addr_w_wire_18;        

  wire [7:0] addr_w_wire_19;        

  wire [7:0] addr_w_wire_20;        

  wire [7:0] addr_w_wire_21;        

  wire [7:0] addr_w_wire_22;        

  wire [7:0] addr_w_wire_23;        

  wire [7:0] addr_w_wire_24;        

  wire [7:0] addr_w_wire_25;        

  wire [7:0] addr_w_wire_26;        

  wire [7:0] addr_w_wire_27;        

  wire [7:0] addr_w_wire_28;        

  wire [7:0] addr_w_wire_29;        

  wire [7:0] addr_w_wire_30;        

  wire [7:0] addr_w_wire_31;        

  wire [7:0] addr_w_wire_32;        

  wire [7:0] addr_w_wire_33;        

  wire [7:0] addr_w_wire_34;        

  wire [7:0] addr_w_wire_35;        

  wire [7:0] addr_w_wire_36;        

  wire [7:0] addr_w_wire_37;        

  wire [7:0] addr_w_wire_38;        

  wire [7:0] addr_w_wire_39;        

  wire [7:0] addr_w_wire_40;        

  wire [7:0] addr_w_wire_41;        

  wire [7:0] addr_w_wire_42;        

  wire [7:0] addr_w_wire_43;        

  wire [7:0] addr_w_wire_44;        

  wire [7:0] addr_w_wire_45;        

  wire [7:0] addr_w_wire_46;        

  wire [7:0] addr_w_wire_47;        

  wire [7:0] addr_w_wire_48;        

  wire [7:0] addr_w_wire_49;        

  wire [7:0] addr_w_wire_50;        

  wire [7:0] addr_w_wire_51;        

  wire [7:0] addr_w_wire_52;        

  wire [7:0] addr_w_wire_53;        

  wire [7:0] addr_w_wire_54;        

  wire [7:0] addr_w_wire_55;        

  wire [7:0] addr_w_wire_56;        

  wire [7:0] addr_w_wire_57;        

  wire [7:0] addr_w_wire_58;        

  wire [7:0] addr_w_wire_59;        

  wire [7:0] addr_w_wire_60;        

  wire [7:0] addr_w_wire_61;        

  wire [7:0] addr_w_wire_62;        

  wire [7:0] addr_w_wire_63;        

  wire [7:0] addr_w_wire_64;        

  wire [7:0] addr_w_wire_65;        

  wire [7:0] addr_w_wire_66;        

  wire [7:0] addr_w_wire_67;        

  wire [7:0] addr_w_wire_68;        

  wire [7:0] addr_w_wire_69;        

  wire [7:0] addr_w_wire_70;        

  wire [7:0] addr_w_wire_71;        

  wire [7:0] addr_w_wire_72;        

  wire [7:0] addr_w_wire_73;        

  wire [7:0] addr_w_wire_74;        

  wire [7:0] addr_w_wire_75;        

  wire [7:0] addr_w_wire_76;        

  wire [7:0] addr_w_wire_77;        

  wire [7:0] addr_w_wire_78;        

  wire [7:0] addr_w_wire_79;        

  wire [7:0] addr_w_wire_80;        

  wire [7:0] addr_w_wire_81;        

  wire [7:0] addr_w_wire_82;        

  wire [7:0] addr_w_wire_83;        

  wire [7:0] addr_w_wire_84;        

  wire [7:0] addr_w_wire_85;        

  wire [7:0] addr_w_wire_86;        

  wire [7:0] addr_w_wire_87;        

  wire [7:0] addr_w_wire_88;        

  wire [7:0] addr_w_wire_89;        

  wire [7:0] addr_w_wire_90;        

  wire [7:0] addr_w_wire_91;        

  wire [7:0] addr_w_wire_92;        

  wire [7:0] addr_w_wire_93;        

  wire [7:0] addr_w_wire_94;        

  wire [7:0] addr_w_wire_95;        

  wire [7:0] addr_w_wire_96;        

  wire [7:0] addr_w_wire_97;        

  wire [7:0] addr_w_wire_98;        

  wire [7:0] addr_w_wire_99;        

  wire [7:0] addr_w_wire_100;        

  wire [7:0] addr_w_wire_101;        

  wire [7:0] addr_w_wire_102;        

  wire [7:0] addr_w_wire_103;        

  wire [7:0] addr_w_wire_104;        

  wire [7:0] addr_w_wire_105;        

  wire [7:0] addr_w_wire_106;        

  wire [7:0] addr_w_wire_107;        

  wire [7:0] addr_w_wire_108;        

  wire [7:0] addr_w_wire_109;        

  wire [7:0] addr_w_wire_110;        

  wire [7:0] addr_w_wire_111;        

  wire [7:0] addr_w_wire_112;        

  wire [7:0] addr_w_wire_113;        

  wire [7:0] addr_w_wire_114;        

  wire [7:0] addr_w_wire_115;        

  wire [7:0] addr_w_wire_116;        

  wire [7:0] addr_w_wire_117;        

  wire [7:0] addr_w_wire_118;        

  wire [7:0] addr_w_wire_119;        

  wire [7:0] addr_w_wire_120;        

  wire [7:0] addr_w_wire_121;        

  wire [7:0] addr_w_wire_122;        

  wire [7:0] addr_w_wire_123;        

  wire [7:0] addr_w_wire_124;        

  wire [7:0] addr_w_wire_125;        

  wire [7:0] addr_w_wire_126;        

  wire [7:0] addr_w_wire_127;        

  wire [7:0] addr_w_wire_128;        

  wire [7:0] addr_w_wire_129;        

  wire [7:0] addr_w_wire_130;        

  wire [7:0] addr_w_wire_131;        

  wire [7:0] addr_w_wire_132;        

  wire [7:0] addr_w_wire_133;        

  wire [7:0] addr_w_wire_134;        

  wire [7:0] addr_w_wire_135;        

  wire [7:0] addr_w_wire_136;        

  wire [7:0] addr_w_wire_137;        

  wire [7:0] addr_w_wire_138;        

  wire [7:0] addr_w_wire_139;        

  wire [7:0] addr_w_wire_140;        

  wire [7:0] addr_w_wire_141;        

  wire [7:0] addr_w_wire_142;        

  wire [7:0] addr_w_wire_143;        

  wire [7:0] addr_w_wire_144;        

  wire [7:0] addr_w_wire_145;        

  wire [7:0] addr_w_wire_146;        

  wire [7:0] addr_w_wire_147;        

  wire [7:0] addr_w_wire_148;        

  wire [7:0] addr_w_wire_149;        

  wire [7:0] addr_w_wire_150;        

  wire [7:0] addr_w_wire_151;        

  wire [7:0] addr_w_wire_152;        

  wire [7:0] addr_w_wire_153;        

  wire [7:0] addr_w_wire_154;        

  wire [7:0] addr_w_wire_155;        

  wire [7:0] addr_w_wire_156;        

  wire [7:0] addr_w_wire_157;        

  wire [7:0] addr_w_wire_158;        

  wire [7:0] addr_w_wire_159;        

  wire [7:0] addr_w_wire_160;        

  wire [7:0] addr_w_wire_161;        

  wire [7:0] addr_w_wire_162;        

  wire [7:0] addr_w_wire_163;        

  wire [7:0] addr_w_wire_164;        

  wire [7:0] addr_w_wire_165;        

  wire [7:0] addr_w_wire_166;        

  wire [7:0] addr_w_wire_167;        

  wire [7:0] addr_w_wire_168;        

  wire [7:0] addr_w_wire_169;        

  wire [7:0] addr_w_wire_170;        

  wire [7:0] addr_w_wire_171;        

  wire [7:0] addr_w_wire_172;        

  wire [7:0] addr_w_wire_173;        

  wire [7:0] addr_w_wire_174;        

  wire [7:0] addr_w_wire_175;        

  wire [7:0] addr_w_wire_176;        

  wire [7:0] addr_w_wire_177;        

  wire [7:0] addr_w_wire_178;        

  wire [7:0] addr_w_wire_179;        

  wire [7:0] addr_w_wire_180;        

  wire [7:0] addr_w_wire_181;        

  wire [7:0] addr_w_wire_182;        

  wire [7:0] addr_w_wire_183;        

  wire [7:0] addr_w_wire_184;        

  wire [7:0] addr_w_wire_185;        

  wire [7:0] addr_w_wire_186;        

  wire [7:0] addr_w_wire_187;        

  wire [7:0] addr_w_wire_188;        

  wire [7:0] addr_w_wire_189;        

  wire [7:0] addr_w_wire_190;        

  wire [7:0] addr_w_wire_191;        

  wire [7:0] addr_w_wire_192;        

  wire [7:0] addr_w_wire_193;        

  wire [7:0] addr_w_wire_194;        

  wire [7:0] addr_w_wire_195;        

  wire [7:0] addr_w_wire_196;        

  wire [7:0] addr_w_wire_197;        

  wire [7:0] addr_w_wire_198;        

  wire [7:0] addr_w_wire_199;        

  wire [7:0] addr_w_wire_200;        

  wire [7:0] addr_w_wire_201;        

  wire [7:0] addr_w_wire_202;        

  wire [7:0] addr_w_wire_203;        

  wire [7:0] addr_w_wire_204;        

  wire [7:0] addr_w_wire_205;        

  wire [7:0] addr_w_wire_206;        

  wire [7:0] addr_w_wire_207;        

  wire [7:0] addr_w_wire_208;        

  wire [7:0] addr_w_wire_209;        

  wire [7:0] addr_w_wire_210;        

  wire [7:0] addr_w_wire_211;        

  wire [7:0] addr_w_wire_212;        

  wire [7:0] addr_w_wire_213;        

  wire [7:0] addr_w_wire_214;        

  wire [7:0] addr_w_wire_215;        

  wire [7:0] addr_w_wire_216;        

  wire [7:0] addr_w_wire_217;        

  wire [7:0] addr_w_wire_218;        

  wire [7:0] addr_w_wire_219;        

  wire [7:0] addr_w_wire_220;        

  wire [7:0] addr_w_wire_221;        

  wire [7:0] addr_w_wire_222;        

  wire [7:0] addr_w_wire_223;        

  wire [7:0] addr_w_wire_224;        

  wire [7:0] addr_w_wire_225;        

  wire [7:0] addr_w_wire_226;        

  wire [7:0] addr_w_wire_227;        

  wire [7:0] addr_w_wire_228;        

  wire [7:0] addr_w_wire_229;        

  wire [7:0] addr_w_wire_230;        

  wire [7:0] addr_w_wire_231;        

  wire [7:0] addr_w_wire_232;        

  wire [7:0] addr_w_wire_233;        

  wire [7:0] addr_w_wire_234;        

  wire [7:0] addr_w_wire_235;        

  wire [7:0] addr_w_wire_236;        

  wire [7:0] addr_w_wire_237;        

  wire [7:0] addr_w_wire_238;        

  wire [7:0] addr_w_wire_239;        

  wire [7:0] addr_w_wire_240;        

  wire [7:0] addr_w_wire_241;        

  wire [7:0] addr_w_wire_242;        

  wire [7:0] addr_w_wire_243;        

  wire [7:0] addr_w_wire_244;        

  wire [7:0] addr_w_wire_245;        

  wire [7:0] addr_w_wire_246;        

  wire [7:0] addr_w_wire_247;        

  wire [7:0] addr_w_wire_248;        

  wire [7:0] addr_w_wire_249;        

  wire [7:0] addr_w_wire_250;        

  wire [7:0] addr_w_wire_251;        

  wire [7:0] addr_w_wire_252;        

  wire [7:0] addr_w_wire_253;        

  wire [7:0] addr_w_wire_254;        

  wire [7:0] addr_w_wire_255;        

  wire [7:0] addr_r_wire_0;        

  assign addr_r_wire_0 = counter_in;        

  mem_addr_ctrl_dp256_per0 addr_gen_inst(.in_start(in_start), .counter_in(counter_in), .wen_out(wen_wire), .out_start(out_start_wire), .mem_addr_out_0(addr_wire_0), .mem_addr_out_1(addr_wire_1), .mem_addr_out_2(addr_wire_2), .mem_addr_out_3(addr_wire_3), .mem_addr_out_4(addr_wire_4), .mem_addr_out_5(addr_wire_5), .mem_addr_out_6(addr_wire_6), .mem_addr_out_7(addr_wire_7), .mem_addr_out_8(addr_wire_8), .mem_addr_out_9(addr_wire_9), .mem_addr_out_10(addr_wire_10), .mem_addr_out_11(addr_wire_11), .mem_addr_out_12(addr_wire_12), .mem_addr_out_13(addr_wire_13), .mem_addr_out_14(addr_wire_14), .mem_addr_out_15(addr_wire_15), .mem_addr_out_16(addr_wire_16), .mem_addr_out_17(addr_wire_17), .mem_addr_out_18(addr_wire_18), .mem_addr_out_19(addr_wire_19), .mem_addr_out_20(addr_wire_20), .mem_addr_out_21(addr_wire_21), .mem_addr_out_22(addr_wire_22), .mem_addr_out_23(addr_wire_23), .mem_addr_out_24(addr_wire_24), .mem_addr_out_25(addr_wire_25), .mem_addr_out_26(addr_wire_26), .mem_addr_out_27(addr_wire_27), .mem_addr_out_28(addr_wire_28), .mem_addr_out_29(addr_wire_29), .mem_addr_out_30(addr_wire_30), .mem_addr_out_31(addr_wire_31), .mem_addr_out_32(addr_wire_32), .mem_addr_out_33(addr_wire_33), .mem_addr_out_34(addr_wire_34), .mem_addr_out_35(addr_wire_35), .mem_addr_out_36(addr_wire_36), .mem_addr_out_37(addr_wire_37), .mem_addr_out_38(addr_wire_38), .mem_addr_out_39(addr_wire_39), .mem_addr_out_40(addr_wire_40), .mem_addr_out_41(addr_wire_41), .mem_addr_out_42(addr_wire_42), .mem_addr_out_43(addr_wire_43), .mem_addr_out_44(addr_wire_44), .mem_addr_out_45(addr_wire_45), .mem_addr_out_46(addr_wire_46), .mem_addr_out_47(addr_wire_47), .mem_addr_out_48(addr_wire_48), .mem_addr_out_49(addr_wire_49), .mem_addr_out_50(addr_wire_50), .mem_addr_out_51(addr_wire_51), .mem_addr_out_52(addr_wire_52), .mem_addr_out_53(addr_wire_53), .mem_addr_out_54(addr_wire_54), .mem_addr_out_55(addr_wire_55), .mem_addr_out_56(addr_wire_56), .mem_addr_out_57(addr_wire_57), .mem_addr_out_58(addr_wire_58), .mem_addr_out_59(addr_wire_59), .mem_addr_out_60(addr_wire_60), .mem_addr_out_61(addr_wire_61), .mem_addr_out_62(addr_wire_62), .mem_addr_out_63(addr_wire_63), .mem_addr_out_64(addr_wire_64), .mem_addr_out_65(addr_wire_65), .mem_addr_out_66(addr_wire_66), .mem_addr_out_67(addr_wire_67), .mem_addr_out_68(addr_wire_68), .mem_addr_out_69(addr_wire_69), .mem_addr_out_70(addr_wire_70), .mem_addr_out_71(addr_wire_71), .mem_addr_out_72(addr_wire_72), .mem_addr_out_73(addr_wire_73), .mem_addr_out_74(addr_wire_74), .mem_addr_out_75(addr_wire_75), .mem_addr_out_76(addr_wire_76), .mem_addr_out_77(addr_wire_77), .mem_addr_out_78(addr_wire_78), .mem_addr_out_79(addr_wire_79), .mem_addr_out_80(addr_wire_80), .mem_addr_out_81(addr_wire_81), .mem_addr_out_82(addr_wire_82), .mem_addr_out_83(addr_wire_83), .mem_addr_out_84(addr_wire_84), .mem_addr_out_85(addr_wire_85), .mem_addr_out_86(addr_wire_86), .mem_addr_out_87(addr_wire_87), .mem_addr_out_88(addr_wire_88), .mem_addr_out_89(addr_wire_89), .mem_addr_out_90(addr_wire_90), .mem_addr_out_91(addr_wire_91), .mem_addr_out_92(addr_wire_92), .mem_addr_out_93(addr_wire_93), .mem_addr_out_94(addr_wire_94), .mem_addr_out_95(addr_wire_95), .mem_addr_out_96(addr_wire_96), .mem_addr_out_97(addr_wire_97), .mem_addr_out_98(addr_wire_98), .mem_addr_out_99(addr_wire_99), .mem_addr_out_100(addr_wire_100), .mem_addr_out_101(addr_wire_101), .mem_addr_out_102(addr_wire_102), .mem_addr_out_103(addr_wire_103), .mem_addr_out_104(addr_wire_104), .mem_addr_out_105(addr_wire_105), .mem_addr_out_106(addr_wire_106), .mem_addr_out_107(addr_wire_107), .mem_addr_out_108(addr_wire_108), .mem_addr_out_109(addr_wire_109), .mem_addr_out_110(addr_wire_110), .mem_addr_out_111(addr_wire_111), .mem_addr_out_112(addr_wire_112), .mem_addr_out_113(addr_wire_113), .mem_addr_out_114(addr_wire_114), .mem_addr_out_115(addr_wire_115), .mem_addr_out_116(addr_wire_116), .mem_addr_out_117(addr_wire_117), .mem_addr_out_118(addr_wire_118), .mem_addr_out_119(addr_wire_119), .mem_addr_out_120(addr_wire_120), .mem_addr_out_121(addr_wire_121), .mem_addr_out_122(addr_wire_122), .mem_addr_out_123(addr_wire_123), .mem_addr_out_124(addr_wire_124), .mem_addr_out_125(addr_wire_125), .mem_addr_out_126(addr_wire_126), .mem_addr_out_127(addr_wire_127), .mem_addr_out_128(addr_wire_128), .mem_addr_out_129(addr_wire_129), .mem_addr_out_130(addr_wire_130), .mem_addr_out_131(addr_wire_131), .mem_addr_out_132(addr_wire_132), .mem_addr_out_133(addr_wire_133), .mem_addr_out_134(addr_wire_134), .mem_addr_out_135(addr_wire_135), .mem_addr_out_136(addr_wire_136), .mem_addr_out_137(addr_wire_137), .mem_addr_out_138(addr_wire_138), .mem_addr_out_139(addr_wire_139), .mem_addr_out_140(addr_wire_140), .mem_addr_out_141(addr_wire_141), .mem_addr_out_142(addr_wire_142), .mem_addr_out_143(addr_wire_143), .mem_addr_out_144(addr_wire_144), .mem_addr_out_145(addr_wire_145), .mem_addr_out_146(addr_wire_146), .mem_addr_out_147(addr_wire_147), .mem_addr_out_148(addr_wire_148), .mem_addr_out_149(addr_wire_149), .mem_addr_out_150(addr_wire_150), .mem_addr_out_151(addr_wire_151), .mem_addr_out_152(addr_wire_152), .mem_addr_out_153(addr_wire_153), .mem_addr_out_154(addr_wire_154), .mem_addr_out_155(addr_wire_155), .mem_addr_out_156(addr_wire_156), .mem_addr_out_157(addr_wire_157), .mem_addr_out_158(addr_wire_158), .mem_addr_out_159(addr_wire_159), .mem_addr_out_160(addr_wire_160), .mem_addr_out_161(addr_wire_161), .mem_addr_out_162(addr_wire_162), .mem_addr_out_163(addr_wire_163), .mem_addr_out_164(addr_wire_164), .mem_addr_out_165(addr_wire_165), .mem_addr_out_166(addr_wire_166), .mem_addr_out_167(addr_wire_167), .mem_addr_out_168(addr_wire_168), .mem_addr_out_169(addr_wire_169), .mem_addr_out_170(addr_wire_170), .mem_addr_out_171(addr_wire_171), .mem_addr_out_172(addr_wire_172), .mem_addr_out_173(addr_wire_173), .mem_addr_out_174(addr_wire_174), .mem_addr_out_175(addr_wire_175), .mem_addr_out_176(addr_wire_176), .mem_addr_out_177(addr_wire_177), .mem_addr_out_178(addr_wire_178), .mem_addr_out_179(addr_wire_179), .mem_addr_out_180(addr_wire_180), .mem_addr_out_181(addr_wire_181), .mem_addr_out_182(addr_wire_182), .mem_addr_out_183(addr_wire_183), .mem_addr_out_184(addr_wire_184), .mem_addr_out_185(addr_wire_185), .mem_addr_out_186(addr_wire_186), .mem_addr_out_187(addr_wire_187), .mem_addr_out_188(addr_wire_188), .mem_addr_out_189(addr_wire_189), .mem_addr_out_190(addr_wire_190), .mem_addr_out_191(addr_wire_191), .mem_addr_out_192(addr_wire_192), .mem_addr_out_193(addr_wire_193), .mem_addr_out_194(addr_wire_194), .mem_addr_out_195(addr_wire_195), .mem_addr_out_196(addr_wire_196), .mem_addr_out_197(addr_wire_197), .mem_addr_out_198(addr_wire_198), .mem_addr_out_199(addr_wire_199), .mem_addr_out_200(addr_wire_200), .mem_addr_out_201(addr_wire_201), .mem_addr_out_202(addr_wire_202), .mem_addr_out_203(addr_wire_203), .mem_addr_out_204(addr_wire_204), .mem_addr_out_205(addr_wire_205), .mem_addr_out_206(addr_wire_206), .mem_addr_out_207(addr_wire_207), .mem_addr_out_208(addr_wire_208), .mem_addr_out_209(addr_wire_209), .mem_addr_out_210(addr_wire_210), .mem_addr_out_211(addr_wire_211), .mem_addr_out_212(addr_wire_212), .mem_addr_out_213(addr_wire_213), .mem_addr_out_214(addr_wire_214), .mem_addr_out_215(addr_wire_215), .mem_addr_out_216(addr_wire_216), .mem_addr_out_217(addr_wire_217), .mem_addr_out_218(addr_wire_218), .mem_addr_out_219(addr_wire_219), .mem_addr_out_220(addr_wire_220), .mem_addr_out_221(addr_wire_221), .mem_addr_out_222(addr_wire_222), .mem_addr_out_223(addr_wire_223), .mem_addr_out_224(addr_wire_224), .mem_addr_out_225(addr_wire_225), .mem_addr_out_226(addr_wire_226), .mem_addr_out_227(addr_wire_227), .mem_addr_out_228(addr_wire_228), .mem_addr_out_229(addr_wire_229), .mem_addr_out_230(addr_wire_230), .mem_addr_out_231(addr_wire_231), .mem_addr_out_232(addr_wire_232), .mem_addr_out_233(addr_wire_233), .mem_addr_out_234(addr_wire_234), .mem_addr_out_235(addr_wire_235), .mem_addr_out_236(addr_wire_236), .mem_addr_out_237(addr_wire_237), .mem_addr_out_238(addr_wire_238), .mem_addr_out_239(addr_wire_239), .mem_addr_out_240(addr_wire_240), .mem_addr_out_241(addr_wire_241), .mem_addr_out_242(addr_wire_242), .mem_addr_out_243(addr_wire_243), .mem_addr_out_244(addr_wire_244), .mem_addr_out_245(addr_wire_245), .mem_addr_out_246(addr_wire_246), .mem_addr_out_247(addr_wire_247), .mem_addr_out_248(addr_wire_248), .mem_addr_out_249(addr_wire_249), .mem_addr_out_250(addr_wire_250), .mem_addr_out_251(addr_wire_251), .mem_addr_out_252(addr_wire_252), .mem_addr_out_253(addr_wire_253), .mem_addr_out_254(addr_wire_254), .mem_addr_out_255(addr_wire_255), .clk(clk), .rst(rst));

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_0(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_0), .din(wire_in[0]), .dout(wire_out[0]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_1(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_1), .din(wire_in[1]), .dout(wire_out[1]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_2(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_2), .din(wire_in[2]), .dout(wire_out[2]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_3(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_3), .din(wire_in[3]), .dout(wire_out[3]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_4(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_4), .din(wire_in[4]), .dout(wire_out[4]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_5(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_5), .din(wire_in[5]), .dout(wire_out[5]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_6(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_6), .din(wire_in[6]), .dout(wire_out[6]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_7(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_7), .din(wire_in[7]), .dout(wire_out[7]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_8(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_8), .din(wire_in[8]), .dout(wire_out[8]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_9(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_9), .din(wire_in[9]), .dout(wire_out[9]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_10(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_10), .din(wire_in[10]), .dout(wire_out[10]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_11(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_11), .din(wire_in[11]), .dout(wire_out[11]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_12(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_12), .din(wire_in[12]), .dout(wire_out[12]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_13(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_13), .din(wire_in[13]), .dout(wire_out[13]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_14(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_14), .din(wire_in[14]), .dout(wire_out[14]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_15(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_15), .din(wire_in[15]), .dout(wire_out[15]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_16(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_16), .din(wire_in[16]), .dout(wire_out[16]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_17(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_17), .din(wire_in[17]), .dout(wire_out[17]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_18(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_18), .din(wire_in[18]), .dout(wire_out[18]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_19(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_19), .din(wire_in[19]), .dout(wire_out[19]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_20(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_20), .din(wire_in[20]), .dout(wire_out[20]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_21(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_21), .din(wire_in[21]), .dout(wire_out[21]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_22(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_22), .din(wire_in[22]), .dout(wire_out[22]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_23(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_23), .din(wire_in[23]), .dout(wire_out[23]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_24(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_24), .din(wire_in[24]), .dout(wire_out[24]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_25(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_25), .din(wire_in[25]), .dout(wire_out[25]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_26(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_26), .din(wire_in[26]), .dout(wire_out[26]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_27(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_27), .din(wire_in[27]), .dout(wire_out[27]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_28(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_28), .din(wire_in[28]), .dout(wire_out[28]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_29(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_29), .din(wire_in[29]), .dout(wire_out[29]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_30(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_30), .din(wire_in[30]), .dout(wire_out[30]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_31(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_31), .din(wire_in[31]), .dout(wire_out[31]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_32(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_32), .din(wire_in[32]), .dout(wire_out[32]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_33(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_33), .din(wire_in[33]), .dout(wire_out[33]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_34(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_34), .din(wire_in[34]), .dout(wire_out[34]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_35(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_35), .din(wire_in[35]), .dout(wire_out[35]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_36(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_36), .din(wire_in[36]), .dout(wire_out[36]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_37(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_37), .din(wire_in[37]), .dout(wire_out[37]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_38(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_38), .din(wire_in[38]), .dout(wire_out[38]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_39(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_39), .din(wire_in[39]), .dout(wire_out[39]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_40(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_40), .din(wire_in[40]), .dout(wire_out[40]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_41(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_41), .din(wire_in[41]), .dout(wire_out[41]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_42(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_42), .din(wire_in[42]), .dout(wire_out[42]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_43(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_43), .din(wire_in[43]), .dout(wire_out[43]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_44(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_44), .din(wire_in[44]), .dout(wire_out[44]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_45(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_45), .din(wire_in[45]), .dout(wire_out[45]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_46(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_46), .din(wire_in[46]), .dout(wire_out[46]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_47(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_47), .din(wire_in[47]), .dout(wire_out[47]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_48(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_48), .din(wire_in[48]), .dout(wire_out[48]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_49(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_49), .din(wire_in[49]), .dout(wire_out[49]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_50(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_50), .din(wire_in[50]), .dout(wire_out[50]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_51(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_51), .din(wire_in[51]), .dout(wire_out[51]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_52(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_52), .din(wire_in[52]), .dout(wire_out[52]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_53(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_53), .din(wire_in[53]), .dout(wire_out[53]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_54(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_54), .din(wire_in[54]), .dout(wire_out[54]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_55(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_55), .din(wire_in[55]), .dout(wire_out[55]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_56(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_56), .din(wire_in[56]), .dout(wire_out[56]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_57(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_57), .din(wire_in[57]), .dout(wire_out[57]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_58(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_58), .din(wire_in[58]), .dout(wire_out[58]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_59(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_59), .din(wire_in[59]), .dout(wire_out[59]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_60(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_60), .din(wire_in[60]), .dout(wire_out[60]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_61(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_61), .din(wire_in[61]), .dout(wire_out[61]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_62(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_62), .din(wire_in[62]), .dout(wire_out[62]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_63(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_63), .din(wire_in[63]), .dout(wire_out[63]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_64(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_64), .din(wire_in[64]), .dout(wire_out[64]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_65(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_65), .din(wire_in[65]), .dout(wire_out[65]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_66(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_66), .din(wire_in[66]), .dout(wire_out[66]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_67(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_67), .din(wire_in[67]), .dout(wire_out[67]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_68(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_68), .din(wire_in[68]), .dout(wire_out[68]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_69(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_69), .din(wire_in[69]), .dout(wire_out[69]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_70(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_70), .din(wire_in[70]), .dout(wire_out[70]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_71(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_71), .din(wire_in[71]), .dout(wire_out[71]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_72(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_72), .din(wire_in[72]), .dout(wire_out[72]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_73(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_73), .din(wire_in[73]), .dout(wire_out[73]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_74(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_74), .din(wire_in[74]), .dout(wire_out[74]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_75(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_75), .din(wire_in[75]), .dout(wire_out[75]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_76(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_76), .din(wire_in[76]), .dout(wire_out[76]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_77(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_77), .din(wire_in[77]), .dout(wire_out[77]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_78(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_78), .din(wire_in[78]), .dout(wire_out[78]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_79(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_79), .din(wire_in[79]), .dout(wire_out[79]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_80(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_80), .din(wire_in[80]), .dout(wire_out[80]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_81(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_81), .din(wire_in[81]), .dout(wire_out[81]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_82(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_82), .din(wire_in[82]), .dout(wire_out[82]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_83(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_83), .din(wire_in[83]), .dout(wire_out[83]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_84(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_84), .din(wire_in[84]), .dout(wire_out[84]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_85(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_85), .din(wire_in[85]), .dout(wire_out[85]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_86(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_86), .din(wire_in[86]), .dout(wire_out[86]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_87(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_87), .din(wire_in[87]), .dout(wire_out[87]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_88(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_88), .din(wire_in[88]), .dout(wire_out[88]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_89(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_89), .din(wire_in[89]), .dout(wire_out[89]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_90(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_90), .din(wire_in[90]), .dout(wire_out[90]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_91(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_91), .din(wire_in[91]), .dout(wire_out[91]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_92(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_92), .din(wire_in[92]), .dout(wire_out[92]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_93(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_93), .din(wire_in[93]), .dout(wire_out[93]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_94(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_94), .din(wire_in[94]), .dout(wire_out[94]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_95(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_95), .din(wire_in[95]), .dout(wire_out[95]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_96(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_96), .din(wire_in[96]), .dout(wire_out[96]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_97(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_97), .din(wire_in[97]), .dout(wire_out[97]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_98(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_98), .din(wire_in[98]), .dout(wire_out[98]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_99(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_99), .din(wire_in[99]), .dout(wire_out[99]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_100(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_100), .din(wire_in[100]), .dout(wire_out[100]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_101(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_101), .din(wire_in[101]), .dout(wire_out[101]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_102(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_102), .din(wire_in[102]), .dout(wire_out[102]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_103(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_103), .din(wire_in[103]), .dout(wire_out[103]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_104(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_104), .din(wire_in[104]), .dout(wire_out[104]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_105(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_105), .din(wire_in[105]), .dout(wire_out[105]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_106(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_106), .din(wire_in[106]), .dout(wire_out[106]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_107(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_107), .din(wire_in[107]), .dout(wire_out[107]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_108(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_108), .din(wire_in[108]), .dout(wire_out[108]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_109(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_109), .din(wire_in[109]), .dout(wire_out[109]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_110(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_110), .din(wire_in[110]), .dout(wire_out[110]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_111(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_111), .din(wire_in[111]), .dout(wire_out[111]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_112(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_112), .din(wire_in[112]), .dout(wire_out[112]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_113(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_113), .din(wire_in[113]), .dout(wire_out[113]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_114(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_114), .din(wire_in[114]), .dout(wire_out[114]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_115(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_115), .din(wire_in[115]), .dout(wire_out[115]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_116(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_116), .din(wire_in[116]), .dout(wire_out[116]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_117(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_117), .din(wire_in[117]), .dout(wire_out[117]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_118(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_118), .din(wire_in[118]), .dout(wire_out[118]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_119(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_119), .din(wire_in[119]), .dout(wire_out[119]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_120(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_120), .din(wire_in[120]), .dout(wire_out[120]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_121(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_121), .din(wire_in[121]), .dout(wire_out[121]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_122(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_122), .din(wire_in[122]), .dout(wire_out[122]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_123(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_123), .din(wire_in[123]), .dout(wire_out[123]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_124(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_124), .din(wire_in[124]), .dout(wire_out[124]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_125(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_125), .din(wire_in[125]), .dout(wire_out[125]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_126(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_126), .din(wire_in[126]), .dout(wire_out[126]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_127(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_127), .din(wire_in[127]), .dout(wire_out[127]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_128(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_128), .din(wire_in[128]), .dout(wire_out[128]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_129(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_129), .din(wire_in[129]), .dout(wire_out[129]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_130(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_130), .din(wire_in[130]), .dout(wire_out[130]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_131(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_131), .din(wire_in[131]), .dout(wire_out[131]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_132(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_132), .din(wire_in[132]), .dout(wire_out[132]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_133(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_133), .din(wire_in[133]), .dout(wire_out[133]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_134(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_134), .din(wire_in[134]), .dout(wire_out[134]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_135(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_135), .din(wire_in[135]), .dout(wire_out[135]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_136(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_136), .din(wire_in[136]), .dout(wire_out[136]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_137(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_137), .din(wire_in[137]), .dout(wire_out[137]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_138(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_138), .din(wire_in[138]), .dout(wire_out[138]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_139(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_139), .din(wire_in[139]), .dout(wire_out[139]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_140(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_140), .din(wire_in[140]), .dout(wire_out[140]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_141(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_141), .din(wire_in[141]), .dout(wire_out[141]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_142(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_142), .din(wire_in[142]), .dout(wire_out[142]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_143(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_143), .din(wire_in[143]), .dout(wire_out[143]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_144(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_144), .din(wire_in[144]), .dout(wire_out[144]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_145(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_145), .din(wire_in[145]), .dout(wire_out[145]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_146(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_146), .din(wire_in[146]), .dout(wire_out[146]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_147(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_147), .din(wire_in[147]), .dout(wire_out[147]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_148(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_148), .din(wire_in[148]), .dout(wire_out[148]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_149(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_149), .din(wire_in[149]), .dout(wire_out[149]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_150(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_150), .din(wire_in[150]), .dout(wire_out[150]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_151(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_151), .din(wire_in[151]), .dout(wire_out[151]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_152(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_152), .din(wire_in[152]), .dout(wire_out[152]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_153(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_153), .din(wire_in[153]), .dout(wire_out[153]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_154(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_154), .din(wire_in[154]), .dout(wire_out[154]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_155(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_155), .din(wire_in[155]), .dout(wire_out[155]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_156(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_156), .din(wire_in[156]), .dout(wire_out[156]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_157(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_157), .din(wire_in[157]), .dout(wire_out[157]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_158(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_158), .din(wire_in[158]), .dout(wire_out[158]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_159(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_159), .din(wire_in[159]), .dout(wire_out[159]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_160(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_160), .din(wire_in[160]), .dout(wire_out[160]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_161(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_161), .din(wire_in[161]), .dout(wire_out[161]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_162(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_162), .din(wire_in[162]), .dout(wire_out[162]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_163(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_163), .din(wire_in[163]), .dout(wire_out[163]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_164(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_164), .din(wire_in[164]), .dout(wire_out[164]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_165(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_165), .din(wire_in[165]), .dout(wire_out[165]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_166(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_166), .din(wire_in[166]), .dout(wire_out[166]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_167(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_167), .din(wire_in[167]), .dout(wire_out[167]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_168(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_168), .din(wire_in[168]), .dout(wire_out[168]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_169(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_169), .din(wire_in[169]), .dout(wire_out[169]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_170(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_170), .din(wire_in[170]), .dout(wire_out[170]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_171(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_171), .din(wire_in[171]), .dout(wire_out[171]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_172(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_172), .din(wire_in[172]), .dout(wire_out[172]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_173(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_173), .din(wire_in[173]), .dout(wire_out[173]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_174(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_174), .din(wire_in[174]), .dout(wire_out[174]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_175(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_175), .din(wire_in[175]), .dout(wire_out[175]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_176(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_176), .din(wire_in[176]), .dout(wire_out[176]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_177(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_177), .din(wire_in[177]), .dout(wire_out[177]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_178(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_178), .din(wire_in[178]), .dout(wire_out[178]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_179(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_179), .din(wire_in[179]), .dout(wire_out[179]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_180(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_180), .din(wire_in[180]), .dout(wire_out[180]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_181(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_181), .din(wire_in[181]), .dout(wire_out[181]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_182(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_182), .din(wire_in[182]), .dout(wire_out[182]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_183(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_183), .din(wire_in[183]), .dout(wire_out[183]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_184(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_184), .din(wire_in[184]), .dout(wire_out[184]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_185(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_185), .din(wire_in[185]), .dout(wire_out[185]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_186(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_186), .din(wire_in[186]), .dout(wire_out[186]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_187(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_187), .din(wire_in[187]), .dout(wire_out[187]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_188(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_188), .din(wire_in[188]), .dout(wire_out[188]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_189(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_189), .din(wire_in[189]), .dout(wire_out[189]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_190(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_190), .din(wire_in[190]), .dout(wire_out[190]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_191(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_191), .din(wire_in[191]), .dout(wire_out[191]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_192(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_192), .din(wire_in[192]), .dout(wire_out[192]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_193(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_193), .din(wire_in[193]), .dout(wire_out[193]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_194(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_194), .din(wire_in[194]), .dout(wire_out[194]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_195(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_195), .din(wire_in[195]), .dout(wire_out[195]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_196(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_196), .din(wire_in[196]), .dout(wire_out[196]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_197(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_197), .din(wire_in[197]), .dout(wire_out[197]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_198(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_198), .din(wire_in[198]), .dout(wire_out[198]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_199(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_199), .din(wire_in[199]), .dout(wire_out[199]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_200(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_200), .din(wire_in[200]), .dout(wire_out[200]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_201(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_201), .din(wire_in[201]), .dout(wire_out[201]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_202(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_202), .din(wire_in[202]), .dout(wire_out[202]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_203(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_203), .din(wire_in[203]), .dout(wire_out[203]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_204(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_204), .din(wire_in[204]), .dout(wire_out[204]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_205(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_205), .din(wire_in[205]), .dout(wire_out[205]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_206(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_206), .din(wire_in[206]), .dout(wire_out[206]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_207(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_207), .din(wire_in[207]), .dout(wire_out[207]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_208(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_208), .din(wire_in[208]), .dout(wire_out[208]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_209(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_209), .din(wire_in[209]), .dout(wire_out[209]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_210(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_210), .din(wire_in[210]), .dout(wire_out[210]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_211(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_211), .din(wire_in[211]), .dout(wire_out[211]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_212(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_212), .din(wire_in[212]), .dout(wire_out[212]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_213(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_213), .din(wire_in[213]), .dout(wire_out[213]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_214(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_214), .din(wire_in[214]), .dout(wire_out[214]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_215(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_215), .din(wire_in[215]), .dout(wire_out[215]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_216(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_216), .din(wire_in[216]), .dout(wire_out[216]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_217(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_217), .din(wire_in[217]), .dout(wire_out[217]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_218(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_218), .din(wire_in[218]), .dout(wire_out[218]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_219(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_219), .din(wire_in[219]), .dout(wire_out[219]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_220(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_220), .din(wire_in[220]), .dout(wire_out[220]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_221(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_221), .din(wire_in[221]), .dout(wire_out[221]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_222(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_222), .din(wire_in[222]), .dout(wire_out[222]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_223(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_223), .din(wire_in[223]), .dout(wire_out[223]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_224(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_224), .din(wire_in[224]), .dout(wire_out[224]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_225(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_225), .din(wire_in[225]), .dout(wire_out[225]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_226(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_226), .din(wire_in[226]), .dout(wire_out[226]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_227(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_227), .din(wire_in[227]), .dout(wire_out[227]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_228(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_228), .din(wire_in[228]), .dout(wire_out[228]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_229(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_229), .din(wire_in[229]), .dout(wire_out[229]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_230(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_230), .din(wire_in[230]), .dout(wire_out[230]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_231(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_231), .din(wire_in[231]), .dout(wire_out[231]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_232(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_232), .din(wire_in[232]), .dout(wire_out[232]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_233(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_233), .din(wire_in[233]), .dout(wire_out[233]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_234(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_234), .din(wire_in[234]), .dout(wire_out[234]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_235(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_235), .din(wire_in[235]), .dout(wire_out[235]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_236(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_236), .din(wire_in[236]), .dout(wire_out[236]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_237(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_237), .din(wire_in[237]), .dout(wire_out[237]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_238(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_238), .din(wire_in[238]), .dout(wire_out[238]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_239(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_239), .din(wire_in[239]), .dout(wire_out[239]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_240(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_240), .din(wire_in[240]), .dout(wire_out[240]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_241(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_241), .din(wire_in[241]), .dout(wire_out[241]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_242(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_242), .din(wire_in[242]), .dout(wire_out[242]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_243(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_243), .din(wire_in[243]), .dout(wire_out[243]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_244(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_244), .din(wire_in[244]), .dout(wire_out[244]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_245(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_245), .din(wire_in[245]), .dout(wire_out[245]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_246(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_246), .din(wire_in[246]), .dout(wire_out[246]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_247(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_247), .din(wire_in[247]), .dout(wire_out[247]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_248(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_248), .din(wire_in[248]), .dout(wire_out[248]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_249(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_249), .din(wire_in[249]), .dout(wire_out[249]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_250(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_250), .din(wire_in[250]), .dout(wire_out[250]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_251(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_251), .din(wire_in[251]), .dout(wire_out[251]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_252(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_252), .din(wire_in[252]), .dout(wire_out[252]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_253(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_253), .din(wire_in[253]), .dout(wire_out[253]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_254(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_254), .din(wire_in[254]), .dout(wire_out[254]), .clk(clk) );

  dist_ram_dp #(.DATA_WIDTH(0), .ADDR_WIDTH(8)) 
         ram_inst_255(.wen(wen_wire), .addr_r(addr_r_wire_0), .addr_w(addr_w_wire_255), .din(wire_in[255]), .dout(wire_out[255]), .clk(clk) );

  
  always@(posedge clk)             
  begin                            
    if(rst) begin                    
      outData_0 <= 0;    
      outData_1 <= 0;    
      outData_2 <= 0;    
      outData_3 <= 0;    
      outData_4 <= 0;    
      outData_5 <= 0;    
      outData_6 <= 0;    
      outData_7 <= 0;    
      outData_8 <= 0;    
      outData_9 <= 0;    
      outData_10 <= 0;    
      outData_11 <= 0;    
      outData_12 <= 0;    
      outData_13 <= 0;    
      outData_14 <= 0;    
      outData_15 <= 0;    
      outData_16 <= 0;    
      outData_17 <= 0;    
      outData_18 <= 0;    
      outData_19 <= 0;    
      outData_20 <= 0;    
      outData_21 <= 0;    
      outData_22 <= 0;    
      outData_23 <= 0;    
      outData_24 <= 0;    
      outData_25 <= 0;    
      outData_26 <= 0;    
      outData_27 <= 0;    
      outData_28 <= 0;    
      outData_29 <= 0;    
      outData_30 <= 0;    
      outData_31 <= 0;    
      outData_32 <= 0;    
      outData_33 <= 0;    
      outData_34 <= 0;    
      outData_35 <= 0;    
      outData_36 <= 0;    
      outData_37 <= 0;    
      outData_38 <= 0;    
      outData_39 <= 0;    
      outData_40 <= 0;    
      outData_41 <= 0;    
      outData_42 <= 0;    
      outData_43 <= 0;    
      outData_44 <= 0;    
      outData_45 <= 0;    
      outData_46 <= 0;    
      outData_47 <= 0;    
      outData_48 <= 0;    
      outData_49 <= 0;    
      outData_50 <= 0;    
      outData_51 <= 0;    
      outData_52 <= 0;    
      outData_53 <= 0;    
      outData_54 <= 0;    
      outData_55 <= 0;    
      outData_56 <= 0;    
      outData_57 <= 0;    
      outData_58 <= 0;    
      outData_59 <= 0;    
      outData_60 <= 0;    
      outData_61 <= 0;    
      outData_62 <= 0;    
      outData_63 <= 0;    
      outData_64 <= 0;    
      outData_65 <= 0;    
      outData_66 <= 0;    
      outData_67 <= 0;    
      outData_68 <= 0;    
      outData_69 <= 0;    
      outData_70 <= 0;    
      outData_71 <= 0;    
      outData_72 <= 0;    
      outData_73 <= 0;    
      outData_74 <= 0;    
      outData_75 <= 0;    
      outData_76 <= 0;    
      outData_77 <= 0;    
      outData_78 <= 0;    
      outData_79 <= 0;    
      outData_80 <= 0;    
      outData_81 <= 0;    
      outData_82 <= 0;    
      outData_83 <= 0;    
      outData_84 <= 0;    
      outData_85 <= 0;    
      outData_86 <= 0;    
      outData_87 <= 0;    
      outData_88 <= 0;    
      outData_89 <= 0;    
      outData_90 <= 0;    
      outData_91 <= 0;    
      outData_92 <= 0;    
      outData_93 <= 0;    
      outData_94 <= 0;    
      outData_95 <= 0;    
      outData_96 <= 0;    
      outData_97 <= 0;    
      outData_98 <= 0;    
      outData_99 <= 0;    
      outData_100 <= 0;    
      outData_101 <= 0;    
      outData_102 <= 0;    
      outData_103 <= 0;    
      outData_104 <= 0;    
      outData_105 <= 0;    
      outData_106 <= 0;    
      outData_107 <= 0;    
      outData_108 <= 0;    
      outData_109 <= 0;    
      outData_110 <= 0;    
      outData_111 <= 0;    
      outData_112 <= 0;    
      outData_113 <= 0;    
      outData_114 <= 0;    
      outData_115 <= 0;    
      outData_116 <= 0;    
      outData_117 <= 0;    
      outData_118 <= 0;    
      outData_119 <= 0;    
      outData_120 <= 0;    
      outData_121 <= 0;    
      outData_122 <= 0;    
      outData_123 <= 0;    
      outData_124 <= 0;    
      outData_125 <= 0;    
      outData_126 <= 0;    
      outData_127 <= 0;    
      outData_128 <= 0;    
      outData_129 <= 0;    
      outData_130 <= 0;    
      outData_131 <= 0;    
      outData_132 <= 0;    
      outData_133 <= 0;    
      outData_134 <= 0;    
      outData_135 <= 0;    
      outData_136 <= 0;    
      outData_137 <= 0;    
      outData_138 <= 0;    
      outData_139 <= 0;    
      outData_140 <= 0;    
      outData_141 <= 0;    
      outData_142 <= 0;    
      outData_143 <= 0;    
      outData_144 <= 0;    
      outData_145 <= 0;    
      outData_146 <= 0;    
      outData_147 <= 0;    
      outData_148 <= 0;    
      outData_149 <= 0;    
      outData_150 <= 0;    
      outData_151 <= 0;    
      outData_152 <= 0;    
      outData_153 <= 0;    
      outData_154 <= 0;    
      outData_155 <= 0;    
      outData_156 <= 0;    
      outData_157 <= 0;    
      outData_158 <= 0;    
      outData_159 <= 0;    
      outData_160 <= 0;    
      outData_161 <= 0;    
      outData_162 <= 0;    
      outData_163 <= 0;    
      outData_164 <= 0;    
      outData_165 <= 0;    
      outData_166 <= 0;    
      outData_167 <= 0;    
      outData_168 <= 0;    
      outData_169 <= 0;    
      outData_170 <= 0;    
      outData_171 <= 0;    
      outData_172 <= 0;    
      outData_173 <= 0;    
      outData_174 <= 0;    
      outData_175 <= 0;    
      outData_176 <= 0;    
      outData_177 <= 0;    
      outData_178 <= 0;    
      outData_179 <= 0;    
      outData_180 <= 0;    
      outData_181 <= 0;    
      outData_182 <= 0;    
      outData_183 <= 0;    
      outData_184 <= 0;    
      outData_185 <= 0;    
      outData_186 <= 0;    
      outData_187 <= 0;    
      outData_188 <= 0;    
      outData_189 <= 0;    
      outData_190 <= 0;    
      outData_191 <= 0;    
      outData_192 <= 0;    
      outData_193 <= 0;    
      outData_194 <= 0;    
      outData_195 <= 0;    
      outData_196 <= 0;    
      outData_197 <= 0;    
      outData_198 <= 0;    
      outData_199 <= 0;    
      outData_200 <= 0;    
      outData_201 <= 0;    
      outData_202 <= 0;    
      outData_203 <= 0;    
      outData_204 <= 0;    
      outData_205 <= 0;    
      outData_206 <= 0;    
      outData_207 <= 0;    
      outData_208 <= 0;    
      outData_209 <= 0;    
      outData_210 <= 0;    
      outData_211 <= 0;    
      outData_212 <= 0;    
      outData_213 <= 0;    
      outData_214 <= 0;    
      outData_215 <= 0;    
      outData_216 <= 0;    
      outData_217 <= 0;    
      outData_218 <= 0;    
      outData_219 <= 0;    
      outData_220 <= 0;    
      outData_221 <= 0;    
      outData_222 <= 0;    
      outData_223 <= 0;    
      outData_224 <= 0;    
      outData_225 <= 0;    
      outData_226 <= 0;    
      outData_227 <= 0;    
      outData_228 <= 0;    
      outData_229 <= 0;    
      outData_230 <= 0;    
      outData_231 <= 0;    
      outData_232 <= 0;    
      outData_233 <= 0;    
      outData_234 <= 0;    
      outData_235 <= 0;    
      outData_236 <= 0;    
      outData_237 <= 0;    
      outData_238 <= 0;    
      outData_239 <= 0;    
      outData_240 <= 0;    
      outData_241 <= 0;    
      outData_242 <= 0;    
      outData_243 <= 0;    
      outData_244 <= 0;    
      outData_245 <= 0;    
      outData_246 <= 0;    
      outData_247 <= 0;    
      outData_248 <= 0;    
      outData_249 <= 0;    
      outData_250 <= 0;    
      outData_251 <= 0;    
      outData_252 <= 0;    
      outData_253 <= 0;    
      outData_254 <= 0;    
      outData_255 <= 0;    
      out_start <= 1'b0;              
      end
    else begin                        
      outData_0 <= wire_out[0];    
      outData_1 <= wire_out[1];    
      outData_2 <= wire_out[2];    
      outData_3 <= wire_out[3];    
      outData_4 <= wire_out[4];    
      outData_5 <= wire_out[5];    
      outData_6 <= wire_out[6];    
      outData_7 <= wire_out[7];    
      outData_8 <= wire_out[8];    
      outData_9 <= wire_out[9];    
      outData_10 <= wire_out[10];    
      outData_11 <= wire_out[11];    
      outData_12 <= wire_out[12];    
      outData_13 <= wire_out[13];    
      outData_14 <= wire_out[14];    
      outData_15 <= wire_out[15];    
      outData_16 <= wire_out[16];    
      outData_17 <= wire_out[17];    
      outData_18 <= wire_out[18];    
      outData_19 <= wire_out[19];    
      outData_20 <= wire_out[20];    
      outData_21 <= wire_out[21];    
      outData_22 <= wire_out[22];    
      outData_23 <= wire_out[23];    
      outData_24 <= wire_out[24];    
      outData_25 <= wire_out[25];    
      outData_26 <= wire_out[26];    
      outData_27 <= wire_out[27];    
      outData_28 <= wire_out[28];    
      outData_29 <= wire_out[29];    
      outData_30 <= wire_out[30];    
      outData_31 <= wire_out[31];    
      outData_32 <= wire_out[32];    
      outData_33 <= wire_out[33];    
      outData_34 <= wire_out[34];    
      outData_35 <= wire_out[35];    
      outData_36 <= wire_out[36];    
      outData_37 <= wire_out[37];    
      outData_38 <= wire_out[38];    
      outData_39 <= wire_out[39];    
      outData_40 <= wire_out[40];    
      outData_41 <= wire_out[41];    
      outData_42 <= wire_out[42];    
      outData_43 <= wire_out[43];    
      outData_44 <= wire_out[44];    
      outData_45 <= wire_out[45];    
      outData_46 <= wire_out[46];    
      outData_47 <= wire_out[47];    
      outData_48 <= wire_out[48];    
      outData_49 <= wire_out[49];    
      outData_50 <= wire_out[50];    
      outData_51 <= wire_out[51];    
      outData_52 <= wire_out[52];    
      outData_53 <= wire_out[53];    
      outData_54 <= wire_out[54];    
      outData_55 <= wire_out[55];    
      outData_56 <= wire_out[56];    
      outData_57 <= wire_out[57];    
      outData_58 <= wire_out[58];    
      outData_59 <= wire_out[59];    
      outData_60 <= wire_out[60];    
      outData_61 <= wire_out[61];    
      outData_62 <= wire_out[62];    
      outData_63 <= wire_out[63];    
      outData_64 <= wire_out[64];    
      outData_65 <= wire_out[65];    
      outData_66 <= wire_out[66];    
      outData_67 <= wire_out[67];    
      outData_68 <= wire_out[68];    
      outData_69 <= wire_out[69];    
      outData_70 <= wire_out[70];    
      outData_71 <= wire_out[71];    
      outData_72 <= wire_out[72];    
      outData_73 <= wire_out[73];    
      outData_74 <= wire_out[74];    
      outData_75 <= wire_out[75];    
      outData_76 <= wire_out[76];    
      outData_77 <= wire_out[77];    
      outData_78 <= wire_out[78];    
      outData_79 <= wire_out[79];    
      outData_80 <= wire_out[80];    
      outData_81 <= wire_out[81];    
      outData_82 <= wire_out[82];    
      outData_83 <= wire_out[83];    
      outData_84 <= wire_out[84];    
      outData_85 <= wire_out[85];    
      outData_86 <= wire_out[86];    
      outData_87 <= wire_out[87];    
      outData_88 <= wire_out[88];    
      outData_89 <= wire_out[89];    
      outData_90 <= wire_out[90];    
      outData_91 <= wire_out[91];    
      outData_92 <= wire_out[92];    
      outData_93 <= wire_out[93];    
      outData_94 <= wire_out[94];    
      outData_95 <= wire_out[95];    
      outData_96 <= wire_out[96];    
      outData_97 <= wire_out[97];    
      outData_98 <= wire_out[98];    
      outData_99 <= wire_out[99];    
      outData_100 <= wire_out[100];    
      outData_101 <= wire_out[101];    
      outData_102 <= wire_out[102];    
      outData_103 <= wire_out[103];    
      outData_104 <= wire_out[104];    
      outData_105 <= wire_out[105];    
      outData_106 <= wire_out[106];    
      outData_107 <= wire_out[107];    
      outData_108 <= wire_out[108];    
      outData_109 <= wire_out[109];    
      outData_110 <= wire_out[110];    
      outData_111 <= wire_out[111];    
      outData_112 <= wire_out[112];    
      outData_113 <= wire_out[113];    
      outData_114 <= wire_out[114];    
      outData_115 <= wire_out[115];    
      outData_116 <= wire_out[116];    
      outData_117 <= wire_out[117];    
      outData_118 <= wire_out[118];    
      outData_119 <= wire_out[119];    
      outData_120 <= wire_out[120];    
      outData_121 <= wire_out[121];    
      outData_122 <= wire_out[122];    
      outData_123 <= wire_out[123];    
      outData_124 <= wire_out[124];    
      outData_125 <= wire_out[125];    
      outData_126 <= wire_out[126];    
      outData_127 <= wire_out[127];    
      outData_128 <= wire_out[128];    
      outData_129 <= wire_out[129];    
      outData_130 <= wire_out[130];    
      outData_131 <= wire_out[131];    
      outData_132 <= wire_out[132];    
      outData_133 <= wire_out[133];    
      outData_134 <= wire_out[134];    
      outData_135 <= wire_out[135];    
      outData_136 <= wire_out[136];    
      outData_137 <= wire_out[137];    
      outData_138 <= wire_out[138];    
      outData_139 <= wire_out[139];    
      outData_140 <= wire_out[140];    
      outData_141 <= wire_out[141];    
      outData_142 <= wire_out[142];    
      outData_143 <= wire_out[143];    
      outData_144 <= wire_out[144];    
      outData_145 <= wire_out[145];    
      outData_146 <= wire_out[146];    
      outData_147 <= wire_out[147];    
      outData_148 <= wire_out[148];    
      outData_149 <= wire_out[149];    
      outData_150 <= wire_out[150];    
      outData_151 <= wire_out[151];    
      outData_152 <= wire_out[152];    
      outData_153 <= wire_out[153];    
      outData_154 <= wire_out[154];    
      outData_155 <= wire_out[155];    
      outData_156 <= wire_out[156];    
      outData_157 <= wire_out[157];    
      outData_158 <= wire_out[158];    
      outData_159 <= wire_out[159];    
      outData_160 <= wire_out[160];    
      outData_161 <= wire_out[161];    
      outData_162 <= wire_out[162];    
      outData_163 <= wire_out[163];    
      outData_164 <= wire_out[164];    
      outData_165 <= wire_out[165];    
      outData_166 <= wire_out[166];    
      outData_167 <= wire_out[167];    
      outData_168 <= wire_out[168];    
      outData_169 <= wire_out[169];    
      outData_170 <= wire_out[170];    
      outData_171 <= wire_out[171];    
      outData_172 <= wire_out[172];    
      outData_173 <= wire_out[173];    
      outData_174 <= wire_out[174];    
      outData_175 <= wire_out[175];    
      outData_176 <= wire_out[176];    
      outData_177 <= wire_out[177];    
      outData_178 <= wire_out[178];    
      outData_179 <= wire_out[179];    
      outData_180 <= wire_out[180];    
      outData_181 <= wire_out[181];    
      outData_182 <= wire_out[182];    
      outData_183 <= wire_out[183];    
      outData_184 <= wire_out[184];    
      outData_185 <= wire_out[185];    
      outData_186 <= wire_out[186];    
      outData_187 <= wire_out[187];    
      outData_188 <= wire_out[188];    
      outData_189 <= wire_out[189];    
      outData_190 <= wire_out[190];    
      outData_191 <= wire_out[191];    
      outData_192 <= wire_out[192];    
      outData_193 <= wire_out[193];    
      outData_194 <= wire_out[194];    
      outData_195 <= wire_out[195];    
      outData_196 <= wire_out[196];    
      outData_197 <= wire_out[197];    
      outData_198 <= wire_out[198];    
      outData_199 <= wire_out[199];    
      outData_200 <= wire_out[200];    
      outData_201 <= wire_out[201];    
      outData_202 <= wire_out[202];    
      outData_203 <= wire_out[203];    
      outData_204 <= wire_out[204];    
      outData_205 <= wire_out[205];    
      outData_206 <= wire_out[206];    
      outData_207 <= wire_out[207];    
      outData_208 <= wire_out[208];    
      outData_209 <= wire_out[209];    
      outData_210 <= wire_out[210];    
      outData_211 <= wire_out[211];    
      outData_212 <= wire_out[212];    
      outData_213 <= wire_out[213];    
      outData_214 <= wire_out[214];    
      outData_215 <= wire_out[215];    
      outData_216 <= wire_out[216];    
      outData_217 <= wire_out[217];    
      outData_218 <= wire_out[218];    
      outData_219 <= wire_out[219];    
      outData_220 <= wire_out[220];    
      outData_221 <= wire_out[221];    
      outData_222 <= wire_out[222];    
      outData_223 <= wire_out[223];    
      outData_224 <= wire_out[224];    
      outData_225 <= wire_out[225];    
      outData_226 <= wire_out[226];    
      outData_227 <= wire_out[227];    
      outData_228 <= wire_out[228];    
      outData_229 <= wire_out[229];    
      outData_230 <= wire_out[230];    
      outData_231 <= wire_out[231];    
      outData_232 <= wire_out[232];    
      outData_233 <= wire_out[233];    
      outData_234 <= wire_out[234];    
      outData_235 <= wire_out[235];    
      outData_236 <= wire_out[236];    
      outData_237 <= wire_out[237];    
      outData_238 <= wire_out[238];    
      outData_239 <= wire_out[239];    
      outData_240 <= wire_out[240];    
      outData_241 <= wire_out[241];    
      outData_242 <= wire_out[242];    
      outData_243 <= wire_out[243];    
      outData_244 <= wire_out[244];    
      outData_245 <= wire_out[245];    
      outData_246 <= wire_out[246];    
      outData_247 <= wire_out[247];    
      outData_248 <= wire_out[248];    
      outData_249 <= wire_out[249];    
      outData_250 <= wire_out[250];    
      outData_251 <= wire_out[251];    
      outData_252 <= wire_out[252];    
      outData_253 <= wire_out[253];    
      outData_254 <= wire_out[254];    
      outData_255 <= wire_out[255];    
      out_start <= out_start_wire;    
      end
  end                              

endmodule                        


module per_dp256_0_r(
inData_0,
inData_1,
inData_2,
inData_3,
inData_4,
inData_5,
inData_6,
inData_7,
inData_8,
inData_9,
inData_10,
inData_11,
inData_12,
inData_13,
inData_14,
inData_15,
inData_16,
inData_17,
inData_18,
inData_19,
inData_20,
inData_21,
inData_22,
inData_23,
inData_24,
inData_25,
inData_26,
inData_27,
inData_28,
inData_29,
inData_30,
inData_31,
inData_32,
inData_33,
inData_34,
inData_35,
inData_36,
inData_37,
inData_38,
inData_39,
inData_40,
inData_41,
inData_42,
inData_43,
inData_44,
inData_45,
inData_46,
inData_47,
inData_48,
inData_49,
inData_50,
inData_51,
inData_52,
inData_53,
inData_54,
inData_55,
inData_56,
inData_57,
inData_58,
inData_59,
inData_60,
inData_61,
inData_62,
inData_63,
inData_64,
inData_65,
inData_66,
inData_67,
inData_68,
inData_69,
inData_70,
inData_71,
inData_72,
inData_73,
inData_74,
inData_75,
inData_76,
inData_77,
inData_78,
inData_79,
inData_80,
inData_81,
inData_82,
inData_83,
inData_84,
inData_85,
inData_86,
inData_87,
inData_88,
inData_89,
inData_90,
inData_91,
inData_92,
inData_93,
inData_94,
inData_95,
inData_96,
inData_97,
inData_98,
inData_99,
inData_100,
inData_101,
inData_102,
inData_103,
inData_104,
inData_105,
inData_106,
inData_107,
inData_108,
inData_109,
inData_110,
inData_111,
inData_112,
inData_113,
inData_114,
inData_115,
inData_116,
inData_117,
inData_118,
inData_119,
inData_120,
inData_121,
inData_122,
inData_123,
inData_124,
inData_125,
inData_126,
inData_127,
inData_128,
inData_129,
inData_130,
inData_131,
inData_132,
inData_133,
inData_134,
inData_135,
inData_136,
inData_137,
inData_138,
inData_139,
inData_140,
inData_141,
inData_142,
inData_143,
inData_144,
inData_145,
inData_146,
inData_147,
inData_148,
inData_149,
inData_150,
inData_151,
inData_152,
inData_153,
inData_154,
inData_155,
inData_156,
inData_157,
inData_158,
inData_159,
inData_160,
inData_161,
inData_162,
inData_163,
inData_164,
inData_165,
inData_166,
inData_167,
inData_168,
inData_169,
inData_170,
inData_171,
inData_172,
inData_173,
inData_174,
inData_175,
inData_176,
inData_177,
inData_178,
inData_179,
inData_180,
inData_181,
inData_182,
inData_183,
inData_184,
inData_185,
inData_186,
inData_187,
inData_188,
inData_189,
inData_190,
inData_191,
inData_192,
inData_193,
inData_194,
inData_195,
inData_196,
inData_197,
inData_198,
inData_199,
inData_200,
inData_201,
inData_202,
inData_203,
inData_204,
inData_205,
inData_206,
inData_207,
inData_208,
inData_209,
inData_210,
inData_211,
inData_212,
inData_213,
inData_214,
inData_215,
inData_216,
inData_217,
inData_218,
inData_219,
inData_220,
inData_221,
inData_222,
inData_223,
inData_224,
inData_225,
inData_226,
inData_227,
inData_228,
inData_229,
inData_230,
inData_231,
inData_232,
inData_233,
inData_234,
inData_235,
inData_236,
inData_237,
inData_238,
inData_239,
inData_240,
inData_241,
inData_242,
inData_243,
inData_244,
inData_245,
inData_246,
inData_247,
inData_248,
inData_249,
inData_250,
inData_251,
inData_252,
inData_253,
inData_254,
inData_255,
outData_0,
outData_1,
outData_2,
outData_3,
outData_4,
outData_5,
outData_6,
outData_7,
outData_8,
outData_9,
outData_10,
outData_11,
outData_12,
outData_13,
outData_14,
outData_15,
outData_16,
outData_17,
outData_18,
outData_19,
outData_20,
outData_21,
outData_22,
outData_23,
outData_24,
outData_25,
outData_26,
outData_27,
outData_28,
outData_29,
outData_30,
outData_31,
outData_32,
outData_33,
outData_34,
outData_35,
outData_36,
outData_37,
outData_38,
outData_39,
outData_40,
outData_41,
outData_42,
outData_43,
outData_44,
outData_45,
outData_46,
outData_47,
outData_48,
outData_49,
outData_50,
outData_51,
outData_52,
outData_53,
outData_54,
outData_55,
outData_56,
outData_57,
outData_58,
outData_59,
outData_60,
outData_61,
outData_62,
outData_63,
outData_64,
outData_65,
outData_66,
outData_67,
outData_68,
outData_69,
outData_70,
outData_71,
outData_72,
outData_73,
outData_74,
outData_75,
outData_76,
outData_77,
outData_78,
outData_79,
outData_80,
outData_81,
outData_82,
outData_83,
outData_84,
outData_85,
outData_86,
outData_87,
outData_88,
outData_89,
outData_90,
outData_91,
outData_92,
outData_93,
outData_94,
outData_95,
outData_96,
outData_97,
outData_98,
outData_99,
outData_100,
outData_101,
outData_102,
outData_103,
outData_104,
outData_105,
outData_106,
outData_107,
outData_108,
outData_109,
outData_110,
outData_111,
outData_112,
outData_113,
outData_114,
outData_115,
outData_116,
outData_117,
outData_118,
outData_119,
outData_120,
outData_121,
outData_122,
outData_123,
outData_124,
outData_125,
outData_126,
outData_127,
outData_128,
outData_129,
outData_130,
outData_131,
outData_132,
outData_133,
outData_134,
outData_135,
outData_136,
outData_137,
outData_138,
outData_139,
outData_140,
outData_141,
outData_142,
outData_143,
outData_144,
outData_145,
outData_146,
outData_147,
outData_148,
outData_149,
outData_150,
outData_151,
outData_152,
outData_153,
outData_154,
outData_155,
outData_156,
outData_157,
outData_158,
outData_159,
outData_160,
outData_161,
outData_162,
outData_163,
outData_164,
outData_165,
outData_166,
outData_167,
outData_168,
outData_169,
outData_170,
outData_171,
outData_172,
outData_173,
outData_174,
outData_175,
outData_176,
outData_177,
outData_178,
outData_179,
outData_180,
outData_181,
outData_182,
outData_183,
outData_184,
outData_185,
outData_186,
outData_187,
outData_188,
outData_189,
outData_190,
outData_191,
outData_192,
outData_193,
outData_194,
outData_195,
outData_196,
outData_197,
outData_198,
outData_199,
outData_200,
outData_201,
outData_202,
outData_203,
outData_204,
outData_205,
outData_206,
outData_207,
outData_208,
outData_209,
outData_210,
outData_211,
outData_212,
outData_213,
outData_214,
outData_215,
outData_216,
outData_217,
outData_218,
outData_219,
outData_220,
outData_221,
outData_222,
outData_223,
outData_224,
outData_225,
outData_226,
outData_227,
outData_228,
outData_229,
outData_230,
outData_231,
outData_232,
outData_233,
outData_234,
outData_235,
outData_236,
outData_237,
outData_238,
outData_239,
outData_240,
outData_241,
outData_242,
outData_243,
outData_244,
outData_245,
outData_246,
outData_247,
outData_248,
outData_249,
outData_250,
outData_251,
outData_252,
outData_253,
outData_254,
outData_255,
in_start,                        
out_start,                       
clk,                             
rst                              
);                               
  parameter DATA_WIDTH = 54;                                
  input in_start, clk, rst;        
  input [DATA_WIDTH-1:0] inData_0,
      inData_1,
      inData_2,
      inData_3,
      inData_4,
      inData_5,
      inData_6,
      inData_7,
      inData_8,
      inData_9,
      inData_10,
      inData_11,
      inData_12,
      inData_13,
      inData_14,
      inData_15,
      inData_16,
      inData_17,
      inData_18,
      inData_19,
      inData_20,
      inData_21,
      inData_22,
      inData_23,
      inData_24,
      inData_25,
      inData_26,
      inData_27,
      inData_28,
      inData_29,
      inData_30,
      inData_31,
      inData_32,
      inData_33,
      inData_34,
      inData_35,
      inData_36,
      inData_37,
      inData_38,
      inData_39,
      inData_40,
      inData_41,
      inData_42,
      inData_43,
      inData_44,
      inData_45,
      inData_46,
      inData_47,
      inData_48,
      inData_49,
      inData_50,
      inData_51,
      inData_52,
      inData_53,
      inData_54,
      inData_55,
      inData_56,
      inData_57,
      inData_58,
      inData_59,
      inData_60,
      inData_61,
      inData_62,
      inData_63,
      inData_64,
      inData_65,
      inData_66,
      inData_67,
      inData_68,
      inData_69,
      inData_70,
      inData_71,
      inData_72,
      inData_73,
      inData_74,
      inData_75,
      inData_76,
      inData_77,
      inData_78,
      inData_79,
      inData_80,
      inData_81,
      inData_82,
      inData_83,
      inData_84,
      inData_85,
      inData_86,
      inData_87,
      inData_88,
      inData_89,
      inData_90,
      inData_91,
      inData_92,
      inData_93,
      inData_94,
      inData_95,
      inData_96,
      inData_97,
      inData_98,
      inData_99,
      inData_100,
      inData_101,
      inData_102,
      inData_103,
      inData_104,
      inData_105,
      inData_106,
      inData_107,
      inData_108,
      inData_109,
      inData_110,
      inData_111,
      inData_112,
      inData_113,
      inData_114,
      inData_115,
      inData_116,
      inData_117,
      inData_118,
      inData_119,
      inData_120,
      inData_121,
      inData_122,
      inData_123,
      inData_124,
      inData_125,
      inData_126,
      inData_127,
      inData_128,
      inData_129,
      inData_130,
      inData_131,
      inData_132,
      inData_133,
      inData_134,
      inData_135,
      inData_136,
      inData_137,
      inData_138,
      inData_139,
      inData_140,
      inData_141,
      inData_142,
      inData_143,
      inData_144,
      inData_145,
      inData_146,
      inData_147,
      inData_148,
      inData_149,
      inData_150,
      inData_151,
      inData_152,
      inData_153,
      inData_154,
      inData_155,
      inData_156,
      inData_157,
      inData_158,
      inData_159,
      inData_160,
      inData_161,
      inData_162,
      inData_163,
      inData_164,
      inData_165,
      inData_166,
      inData_167,
      inData_168,
      inData_169,
      inData_170,
      inData_171,
      inData_172,
      inData_173,
      inData_174,
      inData_175,
      inData_176,
      inData_177,
      inData_178,
      inData_179,
      inData_180,
      inData_181,
      inData_182,
      inData_183,
      inData_184,
      inData_185,
      inData_186,
      inData_187,
      inData_188,
      inData_189,
      inData_190,
      inData_191,
      inData_192,
      inData_193,
      inData_194,
      inData_195,
      inData_196,
      inData_197,
      inData_198,
      inData_199,
      inData_200,
      inData_201,
      inData_202,
      inData_203,
      inData_204,
      inData_205,
      inData_206,
      inData_207,
      inData_208,
      inData_209,
      inData_210,
      inData_211,
      inData_212,
      inData_213,
      inData_214,
      inData_215,
      inData_216,
      inData_217,
      inData_218,
      inData_219,
      inData_220,
      inData_221,
      inData_222,
      inData_223,
      inData_224,
      inData_225,
      inData_226,
      inData_227,
      inData_228,
      inData_229,
      inData_230,
      inData_231,
      inData_232,
      inData_233,
      inData_234,
      inData_235,
      inData_236,
      inData_237,
      inData_238,
      inData_239,
      inData_240,
      inData_241,
      inData_242,
      inData_243,
      inData_244,
      inData_245,
      inData_246,
      inData_247,
      inData_248,
      inData_249,
      inData_250,
      inData_251,
      inData_252,
      inData_253,
      inData_254,
      inData_255;
  output reg [DATA_WIDTH-1:0] outData_0,
      outData_1,
      outData_2,
      outData_3,
      outData_4,
      outData_5,
      outData_6,
      outData_7,
      outData_8,
      outData_9,
      outData_10,
      outData_11,
      outData_12,
      outData_13,
      outData_14,
      outData_15,
      outData_16,
      outData_17,
      outData_18,
      outData_19,
      outData_20,
      outData_21,
      outData_22,
      outData_23,
      outData_24,
      outData_25,
      outData_26,
      outData_27,
      outData_28,
      outData_29,
      outData_30,
      outData_31,
      outData_32,
      outData_33,
      outData_34,
      outData_35,
      outData_36,
      outData_37,
      outData_38,
      outData_39,
      outData_40,
      outData_41,
      outData_42,
      outData_43,
      outData_44,
      outData_45,
      outData_46,
      outData_47,
      outData_48,
      outData_49,
      outData_50,
      outData_51,
      outData_52,
      outData_53,
      outData_54,
      outData_55,
      outData_56,
      outData_57,
      outData_58,
      outData_59,
      outData_60,
      outData_61,
      outData_62,
      outData_63,
      outData_64,
      outData_65,
      outData_66,
      outData_67,
      outData_68,
      outData_69,
      outData_70,
      outData_71,
      outData_72,
      outData_73,
      outData_74,
      outData_75,
      outData_76,
      outData_77,
      outData_78,
      outData_79,
      outData_80,
      outData_81,
      outData_82,
      outData_83,
      outData_84,
      outData_85,
      outData_86,
      outData_87,
      outData_88,
      outData_89,
      outData_90,
      outData_91,
      outData_92,
      outData_93,
      outData_94,
      outData_95,
      outData_96,
      outData_97,
      outData_98,
      outData_99,
      outData_100,
      outData_101,
      outData_102,
      outData_103,
      outData_104,
      outData_105,
      outData_106,
      outData_107,
      outData_108,
      outData_109,
      outData_110,
      outData_111,
      outData_112,
      outData_113,
      outData_114,
      outData_115,
      outData_116,
      outData_117,
      outData_118,
      outData_119,
      outData_120,
      outData_121,
      outData_122,
      outData_123,
      outData_124,
      outData_125,
      outData_126,
      outData_127,
      outData_128,
      outData_129,
      outData_130,
      outData_131,
      outData_132,
      outData_133,
      outData_134,
      outData_135,
      outData_136,
      outData_137,
      outData_138,
      outData_139,
      outData_140,
      outData_141,
      outData_142,
      outData_143,
      outData_144,
      outData_145,
      outData_146,
      outData_147,
      outData_148,
      outData_149,
      outData_150,
      outData_151,
      outData_152,
      outData_153,
      outData_154,
      outData_155,
      outData_156,
      outData_157,
      outData_158,
      outData_159,
      outData_160,
      outData_161,
      outData_162,
      outData_163,
      outData_164,
      outData_165,
      outData_166,
      outData_167,
      outData_168,
      outData_169,
      outData_170,
      outData_171,
      outData_172,
      outData_173,
      outData_174,
      outData_175,
      outData_176,
      outData_177,
      outData_178,
      outData_179,
      outData_180,
      outData_181,
      outData_182,
      outData_183,
      outData_184,
      outData_185,
      outData_186,
      outData_187,
      outData_188,
      outData_189,
      outData_190,
      outData_191,
      outData_192,
      outData_193,
      outData_194,
      outData_195,
      outData_196,
      outData_197,
      outData_198,
      outData_199,
      outData_200,
      outData_201,
      outData_202,
      outData_203,
      outData_204,
      outData_205,
      outData_206,
      outData_207,
      outData_208,
      outData_209,
      outData_210,
      outData_211,
      outData_212,
      outData_213,
      outData_214,
      outData_215,
      outData_216,
      outData_217,
      outData_218,
      outData_219,
      outData_220,
      outData_221,
      outData_222,
      outData_223,
      outData_224,
      outData_225,
      outData_226,
      outData_227,
      outData_228,
      outData_229,
      outData_230,
      outData_231,
      outData_232,
      outData_233,
      outData_234,
      outData_235,
      outData_236,
      outData_237,
      outData_238,
      outData_239,
      outData_240,
      outData_241,
      outData_242,
      outData_243,
      outData_244,
      outData_245,
      outData_246,
      outData_247,
      outData_248,
      outData_249,
      outData_250,
      outData_251,
      outData_252,
      outData_253,
      outData_254,
      outData_255; 
  output reg out_start; 
  
  wire [DATA_WIDTH-1:0] wireIn [255:0];                  
  wire [DATA_WIDTH-1:0] wireOut [255:0];                 
  wire [DATA_WIDTH-1:0] wireOut_LB [255:0];              
  wire [DATA_WIDTH-1:0] wireIn_RB [255:0];               
  wire out_start_LB;               
  wire out_start_MemStage;               
  wire out_start_RB;               

  wire [7:0] counter_out_w;               
  assign wireIn[0] = inData_0;    
  assign wireIn[1] = inData_1;    
  assign wireIn[2] = inData_2;    
  assign wireIn[3] = inData_3;    
  assign wireIn[4] = inData_4;    
  assign wireIn[5] = inData_5;    
  assign wireIn[6] = inData_6;    
  assign wireIn[7] = inData_7;    
  assign wireIn[8] = inData_8;    
  assign wireIn[9] = inData_9;    
  assign wireIn[10] = inData_10;    
  assign wireIn[11] = inData_11;    
  assign wireIn[12] = inData_12;    
  assign wireIn[13] = inData_13;    
  assign wireIn[14] = inData_14;    
  assign wireIn[15] = inData_15;    
  assign wireIn[16] = inData_16;    
  assign wireIn[17] = inData_17;    
  assign wireIn[18] = inData_18;    
  assign wireIn[19] = inData_19;    
  assign wireIn[20] = inData_20;    
  assign wireIn[21] = inData_21;    
  assign wireIn[22] = inData_22;    
  assign wireIn[23] = inData_23;    
  assign wireIn[24] = inData_24;    
  assign wireIn[25] = inData_25;    
  assign wireIn[26] = inData_26;    
  assign wireIn[27] = inData_27;    
  assign wireIn[28] = inData_28;    
  assign wireIn[29] = inData_29;    
  assign wireIn[30] = inData_30;    
  assign wireIn[31] = inData_31;    
  assign wireIn[32] = inData_32;    
  assign wireIn[33] = inData_33;    
  assign wireIn[34] = inData_34;    
  assign wireIn[35] = inData_35;    
  assign wireIn[36] = inData_36;    
  assign wireIn[37] = inData_37;    
  assign wireIn[38] = inData_38;    
  assign wireIn[39] = inData_39;    
  assign wireIn[40] = inData_40;    
  assign wireIn[41] = inData_41;    
  assign wireIn[42] = inData_42;    
  assign wireIn[43] = inData_43;    
  assign wireIn[44] = inData_44;    
  assign wireIn[45] = inData_45;    
  assign wireIn[46] = inData_46;    
  assign wireIn[47] = inData_47;    
  assign wireIn[48] = inData_48;    
  assign wireIn[49] = inData_49;    
  assign wireIn[50] = inData_50;    
  assign wireIn[51] = inData_51;    
  assign wireIn[52] = inData_52;    
  assign wireIn[53] = inData_53;    
  assign wireIn[54] = inData_54;    
  assign wireIn[55] = inData_55;    
  assign wireIn[56] = inData_56;    
  assign wireIn[57] = inData_57;    
  assign wireIn[58] = inData_58;    
  assign wireIn[59] = inData_59;    
  assign wireIn[60] = inData_60;    
  assign wireIn[61] = inData_61;    
  assign wireIn[62] = inData_62;    
  assign wireIn[63] = inData_63;    
  assign wireIn[64] = inData_64;    
  assign wireIn[65] = inData_65;    
  assign wireIn[66] = inData_66;    
  assign wireIn[67] = inData_67;    
  assign wireIn[68] = inData_68;    
  assign wireIn[69] = inData_69;    
  assign wireIn[70] = inData_70;    
  assign wireIn[71] = inData_71;    
  assign wireIn[72] = inData_72;    
  assign wireIn[73] = inData_73;    
  assign wireIn[74] = inData_74;    
  assign wireIn[75] = inData_75;    
  assign wireIn[76] = inData_76;    
  assign wireIn[77] = inData_77;    
  assign wireIn[78] = inData_78;    
  assign wireIn[79] = inData_79;    
  assign wireIn[80] = inData_80;    
  assign wireIn[81] = inData_81;    
  assign wireIn[82] = inData_82;    
  assign wireIn[83] = inData_83;    
  assign wireIn[84] = inData_84;    
  assign wireIn[85] = inData_85;    
  assign wireIn[86] = inData_86;    
  assign wireIn[87] = inData_87;    
  assign wireIn[88] = inData_88;    
  assign wireIn[89] = inData_89;    
  assign wireIn[90] = inData_90;    
  assign wireIn[91] = inData_91;    
  assign wireIn[92] = inData_92;    
  assign wireIn[93] = inData_93;    
  assign wireIn[94] = inData_94;    
  assign wireIn[95] = inData_95;    
  assign wireIn[96] = inData_96;    
  assign wireIn[97] = inData_97;    
  assign wireIn[98] = inData_98;    
  assign wireIn[99] = inData_99;    
  assign wireIn[100] = inData_100;    
  assign wireIn[101] = inData_101;    
  assign wireIn[102] = inData_102;    
  assign wireIn[103] = inData_103;    
  assign wireIn[104] = inData_104;    
  assign wireIn[105] = inData_105;    
  assign wireIn[106] = inData_106;    
  assign wireIn[107] = inData_107;    
  assign wireIn[108] = inData_108;    
  assign wireIn[109] = inData_109;    
  assign wireIn[110] = inData_110;    
  assign wireIn[111] = inData_111;    
  assign wireIn[112] = inData_112;    
  assign wireIn[113] = inData_113;    
  assign wireIn[114] = inData_114;    
  assign wireIn[115] = inData_115;    
  assign wireIn[116] = inData_116;    
  assign wireIn[117] = inData_117;    
  assign wireIn[118] = inData_118;    
  assign wireIn[119] = inData_119;    
  assign wireIn[120] = inData_120;    
  assign wireIn[121] = inData_121;    
  assign wireIn[122] = inData_122;    
  assign wireIn[123] = inData_123;    
  assign wireIn[124] = inData_124;    
  assign wireIn[125] = inData_125;    
  assign wireIn[126] = inData_126;    
  assign wireIn[127] = inData_127;    
  assign wireIn[128] = inData_128;    
  assign wireIn[129] = inData_129;    
  assign wireIn[130] = inData_130;    
  assign wireIn[131] = inData_131;    
  assign wireIn[132] = inData_132;    
  assign wireIn[133] = inData_133;    
  assign wireIn[134] = inData_134;    
  assign wireIn[135] = inData_135;    
  assign wireIn[136] = inData_136;    
  assign wireIn[137] = inData_137;    
  assign wireIn[138] = inData_138;    
  assign wireIn[139] = inData_139;    
  assign wireIn[140] = inData_140;    
  assign wireIn[141] = inData_141;    
  assign wireIn[142] = inData_142;    
  assign wireIn[143] = inData_143;    
  assign wireIn[144] = inData_144;    
  assign wireIn[145] = inData_145;    
  assign wireIn[146] = inData_146;    
  assign wireIn[147] = inData_147;    
  assign wireIn[148] = inData_148;    
  assign wireIn[149] = inData_149;    
  assign wireIn[150] = inData_150;    
  assign wireIn[151] = inData_151;    
  assign wireIn[152] = inData_152;    
  assign wireIn[153] = inData_153;    
  assign wireIn[154] = inData_154;    
  assign wireIn[155] = inData_155;    
  assign wireIn[156] = inData_156;    
  assign wireIn[157] = inData_157;    
  assign wireIn[158] = inData_158;    
  assign wireIn[159] = inData_159;    
  assign wireIn[160] = inData_160;    
  assign wireIn[161] = inData_161;    
  assign wireIn[162] = inData_162;    
  assign wireIn[163] = inData_163;    
  assign wireIn[164] = inData_164;    
  assign wireIn[165] = inData_165;    
  assign wireIn[166] = inData_166;    
  assign wireIn[167] = inData_167;    
  assign wireIn[168] = inData_168;    
  assign wireIn[169] = inData_169;    
  assign wireIn[170] = inData_170;    
  assign wireIn[171] = inData_171;    
  assign wireIn[172] = inData_172;    
  assign wireIn[173] = inData_173;    
  assign wireIn[174] = inData_174;    
  assign wireIn[175] = inData_175;    
  assign wireIn[176] = inData_176;    
  assign wireIn[177] = inData_177;    
  assign wireIn[178] = inData_178;    
  assign wireIn[179] = inData_179;    
  assign wireIn[180] = inData_180;    
  assign wireIn[181] = inData_181;    
  assign wireIn[182] = inData_182;    
  assign wireIn[183] = inData_183;    
  assign wireIn[184] = inData_184;    
  assign wireIn[185] = inData_185;    
  assign wireIn[186] = inData_186;    
  assign wireIn[187] = inData_187;    
  assign wireIn[188] = inData_188;    
  assign wireIn[189] = inData_189;    
  assign wireIn[190] = inData_190;    
  assign wireIn[191] = inData_191;    
  assign wireIn[192] = inData_192;    
  assign wireIn[193] = inData_193;    
  assign wireIn[194] = inData_194;    
  assign wireIn[195] = inData_195;    
  assign wireIn[196] = inData_196;    
  assign wireIn[197] = inData_197;    
  assign wireIn[198] = inData_198;    
  assign wireIn[199] = inData_199;    
  assign wireIn[200] = inData_200;    
  assign wireIn[201] = inData_201;    
  assign wireIn[202] = inData_202;    
  assign wireIn[203] = inData_203;    
  assign wireIn[204] = inData_204;    
  assign wireIn[205] = inData_205;    
  assign wireIn[206] = inData_206;    
  assign wireIn[207] = inData_207;    
  assign wireIn[208] = inData_208;    
  assign wireIn[209] = inData_209;    
  assign wireIn[210] = inData_210;    
  assign wireIn[211] = inData_211;    
  assign wireIn[212] = inData_212;    
  assign wireIn[213] = inData_213;    
  assign wireIn[214] = inData_214;    
  assign wireIn[215] = inData_215;    
  assign wireIn[216] = inData_216;    
  assign wireIn[217] = inData_217;    
  assign wireIn[218] = inData_218;    
  assign wireIn[219] = inData_219;    
  assign wireIn[220] = inData_220;    
  assign wireIn[221] = inData_221;    
  assign wireIn[222] = inData_222;    
  assign wireIn[223] = inData_223;    
  assign wireIn[224] = inData_224;    
  assign wireIn[225] = inData_225;    
  assign wireIn[226] = inData_226;    
  assign wireIn[227] = inData_227;    
  assign wireIn[228] = inData_228;    
  assign wireIn[229] = inData_229;    
  assign wireIn[230] = inData_230;    
  assign wireIn[231] = inData_231;    
  assign wireIn[232] = inData_232;    
  assign wireIn[233] = inData_233;    
  assign wireIn[234] = inData_234;    
  assign wireIn[235] = inData_235;    
  assign wireIn[236] = inData_236;    
  assign wireIn[237] = inData_237;    
  assign wireIn[238] = inData_238;    
  assign wireIn[239] = inData_239;    
  assign wireIn[240] = inData_240;    
  assign wireIn[241] = inData_241;    
  assign wireIn[242] = inData_242;    
  assign wireIn[243] = inData_243;    
  assign wireIn[244] = inData_244;    
  assign wireIn[245] = inData_245;    
  assign wireIn[246] = inData_246;    
  assign wireIn[247] = inData_247;    
  assign wireIn[248] = inData_248;    
  assign wireIn[249] = inData_249;    
  assign wireIn[250] = inData_250;    
  assign wireIn[251] = inData_251;    
  assign wireIn[252] = inData_252;    
  assign wireIn[253] = inData_253;    
  assign wireIn[254] = inData_254;    
  assign wireIn[255] = inData_255;    
  
  counter_512 ctrl_unit(.in_start(in_start), .counter_out(counter_out_w), .clk(clk), .rst(rst));

  ingressStage_p256 ingressStage_p256_inst(.inData_0(wireIn[0]), .inData_1(wireIn[1]), .inData_2(wireIn[2]), .inData_3(wireIn[3]), .inData_4(wireIn[4]), .inData_5(wireIn[5]), .inData_6(wireIn[6]), .inData_7(wireIn[7]), .inData_8(wireIn[8]), .inData_9(wireIn[9]), .inData_10(wireIn[10]), .inData_11(wireIn[11]), .inData_12(wireIn[12]), .inData_13(wireIn[13]), .inData_14(wireIn[14]), .inData_15(wireIn[15]), .inData_16(wireIn[16]), .inData_17(wireIn[17]), .inData_18(wireIn[18]), .inData_19(wireIn[19]), .inData_20(wireIn[20]), .inData_21(wireIn[21]), .inData_22(wireIn[22]), .inData_23(wireIn[23]), .inData_24(wireIn[24]), .inData_25(wireIn[25]), .inData_26(wireIn[26]), .inData_27(wireIn[27]), .inData_28(wireIn[28]), .inData_29(wireIn[29]), .inData_30(wireIn[30]), .inData_31(wireIn[31]), .inData_32(wireIn[32]), .inData_33(wireIn[33]), .inData_34(wireIn[34]), .inData_35(wireIn[35]), .inData_36(wireIn[36]), .inData_37(wireIn[37]), .inData_38(wireIn[38]), .inData_39(wireIn[39]), .inData_40(wireIn[40]), .inData_41(wireIn[41]), .inData_42(wireIn[42]), .inData_43(wireIn[43]), .inData_44(wireIn[44]), .inData_45(wireIn[45]), .inData_46(wireIn[46]), .inData_47(wireIn[47]), .inData_48(wireIn[48]), .inData_49(wireIn[49]), .inData_50(wireIn[50]), .inData_51(wireIn[51]), .inData_52(wireIn[52]), .inData_53(wireIn[53]), .inData_54(wireIn[54]), .inData_55(wireIn[55]), .inData_56(wireIn[56]), .inData_57(wireIn[57]), .inData_58(wireIn[58]), .inData_59(wireIn[59]), .inData_60(wireIn[60]), .inData_61(wireIn[61]), .inData_62(wireIn[62]), .inData_63(wireIn[63]), .inData_64(wireIn[64]), .inData_65(wireIn[65]), .inData_66(wireIn[66]), .inData_67(wireIn[67]), .inData_68(wireIn[68]), .inData_69(wireIn[69]), .inData_70(wireIn[70]), .inData_71(wireIn[71]), .inData_72(wireIn[72]), .inData_73(wireIn[73]), .inData_74(wireIn[74]), .inData_75(wireIn[75]), .inData_76(wireIn[76]), .inData_77(wireIn[77]), .inData_78(wireIn[78]), .inData_79(wireIn[79]), .inData_80(wireIn[80]), .inData_81(wireIn[81]), .inData_82(wireIn[82]), .inData_83(wireIn[83]), .inData_84(wireIn[84]), .inData_85(wireIn[85]), .inData_86(wireIn[86]), .inData_87(wireIn[87]), .inData_88(wireIn[88]), .inData_89(wireIn[89]), .inData_90(wireIn[90]), .inData_91(wireIn[91]), .inData_92(wireIn[92]), .inData_93(wireIn[93]), .inData_94(wireIn[94]), .inData_95(wireIn[95]), .inData_96(wireIn[96]), .inData_97(wireIn[97]), .inData_98(wireIn[98]), .inData_99(wireIn[99]), .inData_100(wireIn[100]), .inData_101(wireIn[101]), .inData_102(wireIn[102]), .inData_103(wireIn[103]), .inData_104(wireIn[104]), .inData_105(wireIn[105]), .inData_106(wireIn[106]), .inData_107(wireIn[107]), .inData_108(wireIn[108]), .inData_109(wireIn[109]), .inData_110(wireIn[110]), .inData_111(wireIn[111]), .inData_112(wireIn[112]), .inData_113(wireIn[113]), .inData_114(wireIn[114]), .inData_115(wireIn[115]), .inData_116(wireIn[116]), .inData_117(wireIn[117]), .inData_118(wireIn[118]), .inData_119(wireIn[119]), .inData_120(wireIn[120]), .inData_121(wireIn[121]), .inData_122(wireIn[122]), .inData_123(wireIn[123]), .inData_124(wireIn[124]), .inData_125(wireIn[125]), .inData_126(wireIn[126]), .inData_127(wireIn[127]), .inData_128(wireIn[128]), .inData_129(wireIn[129]), .inData_130(wireIn[130]), .inData_131(wireIn[131]), .inData_132(wireIn[132]), .inData_133(wireIn[133]), .inData_134(wireIn[134]), .inData_135(wireIn[135]), .inData_136(wireIn[136]), .inData_137(wireIn[137]), .inData_138(wireIn[138]), .inData_139(wireIn[139]), .inData_140(wireIn[140]), .inData_141(wireIn[141]), .inData_142(wireIn[142]), .inData_143(wireIn[143]), .inData_144(wireIn[144]), .inData_145(wireIn[145]), .inData_146(wireIn[146]), .inData_147(wireIn[147]), .inData_148(wireIn[148]), .inData_149(wireIn[149]), .inData_150(wireIn[150]), .inData_151(wireIn[151]), .inData_152(wireIn[152]), .inData_153(wireIn[153]), .inData_154(wireIn[154]), .inData_155(wireIn[155]), .inData_156(wireIn[156]), .inData_157(wireIn[157]), .inData_158(wireIn[158]), .inData_159(wireIn[159]), .inData_160(wireIn[160]), .inData_161(wireIn[161]), .inData_162(wireIn[162]), .inData_163(wireIn[163]), .inData_164(wireIn[164]), .inData_165(wireIn[165]), .inData_166(wireIn[166]), .inData_167(wireIn[167]), .inData_168(wireIn[168]), .inData_169(wireIn[169]), .inData_170(wireIn[170]), .inData_171(wireIn[171]), .inData_172(wireIn[172]), .inData_173(wireIn[173]), .inData_174(wireIn[174]), .inData_175(wireIn[175]), .inData_176(wireIn[176]), .inData_177(wireIn[177]), .inData_178(wireIn[178]), .inData_179(wireIn[179]), .inData_180(wireIn[180]), .inData_181(wireIn[181]), .inData_182(wireIn[182]), .inData_183(wireIn[183]), .inData_184(wireIn[184]), .inData_185(wireIn[185]), .inData_186(wireIn[186]), .inData_187(wireIn[187]), .inData_188(wireIn[188]), .inData_189(wireIn[189]), .inData_190(wireIn[190]), .inData_191(wireIn[191]), .inData_192(wireIn[192]), .inData_193(wireIn[193]), .inData_194(wireIn[194]), .inData_195(wireIn[195]), .inData_196(wireIn[196]), .inData_197(wireIn[197]), .inData_198(wireIn[198]), .inData_199(wireIn[199]), .inData_200(wireIn[200]), .inData_201(wireIn[201]), .inData_202(wireIn[202]), .inData_203(wireIn[203]), .inData_204(wireIn[204]), .inData_205(wireIn[205]), .inData_206(wireIn[206]), .inData_207(wireIn[207]), .inData_208(wireIn[208]), .inData_209(wireIn[209]), .inData_210(wireIn[210]), .inData_211(wireIn[211]), .inData_212(wireIn[212]), .inData_213(wireIn[213]), .inData_214(wireIn[214]), .inData_215(wireIn[215]), .inData_216(wireIn[216]), .inData_217(wireIn[217]), .inData_218(wireIn[218]), .inData_219(wireIn[219]), .inData_220(wireIn[220]), .inData_221(wireIn[221]), .inData_222(wireIn[222]), .inData_223(wireIn[223]), .inData_224(wireIn[224]), .inData_225(wireIn[225]), .inData_226(wireIn[226]), .inData_227(wireIn[227]), .inData_228(wireIn[228]), .inData_229(wireIn[229]), .inData_230(wireIn[230]), .inData_231(wireIn[231]), .inData_232(wireIn[232]), .inData_233(wireIn[233]), .inData_234(wireIn[234]), .inData_235(wireIn[235]), .inData_236(wireIn[236]), .inData_237(wireIn[237]), .inData_238(wireIn[238]), .inData_239(wireIn[239]), .inData_240(wireIn[240]), .inData_241(wireIn[241]), .inData_242(wireIn[242]), .inData_243(wireIn[243]), .inData_244(wireIn[244]), .inData_245(wireIn[245]), .inData_246(wireIn[246]), .inData_247(wireIn[247]), .inData_248(wireIn[248]), .inData_249(wireIn[249]), .inData_250(wireIn[250]), .inData_251(wireIn[251]), .inData_252(wireIn[252]), .inData_253(wireIn[253]), .inData_254(wireIn[254]), .inData_255(wireIn[255]), .outData_0(wireOut_LB[0]), .outData_1(wireOut_LB[1]), .outData_2(wireOut_LB[2]), .outData_3(wireOut_LB[3]), .outData_4(wireOut_LB[4]), .outData_5(wireOut_LB[5]), .outData_6(wireOut_LB[6]), .outData_7(wireOut_LB[7]), .outData_8(wireOut_LB[8]), .outData_9(wireOut_LB[9]), .outData_10(wireOut_LB[10]), .outData_11(wireOut_LB[11]), .outData_12(wireOut_LB[12]), .outData_13(wireOut_LB[13]), .outData_14(wireOut_LB[14]), .outData_15(wireOut_LB[15]), .outData_16(wireOut_LB[16]), .outData_17(wireOut_LB[17]), .outData_18(wireOut_LB[18]), .outData_19(wireOut_LB[19]), .outData_20(wireOut_LB[20]), .outData_21(wireOut_LB[21]), .outData_22(wireOut_LB[22]), .outData_23(wireOut_LB[23]), .outData_24(wireOut_LB[24]), .outData_25(wireOut_LB[25]), .outData_26(wireOut_LB[26]), .outData_27(wireOut_LB[27]), .outData_28(wireOut_LB[28]), .outData_29(wireOut_LB[29]), .outData_30(wireOut_LB[30]), .outData_31(wireOut_LB[31]), .outData_32(wireOut_LB[32]), .outData_33(wireOut_LB[33]), .outData_34(wireOut_LB[34]), .outData_35(wireOut_LB[35]), .outData_36(wireOut_LB[36]), .outData_37(wireOut_LB[37]), .outData_38(wireOut_LB[38]), .outData_39(wireOut_LB[39]), .outData_40(wireOut_LB[40]), .outData_41(wireOut_LB[41]), .outData_42(wireOut_LB[42]), .outData_43(wireOut_LB[43]), .outData_44(wireOut_LB[44]), .outData_45(wireOut_LB[45]), .outData_46(wireOut_LB[46]), .outData_47(wireOut_LB[47]), .outData_48(wireOut_LB[48]), .outData_49(wireOut_LB[49]), .outData_50(wireOut_LB[50]), .outData_51(wireOut_LB[51]), .outData_52(wireOut_LB[52]), .outData_53(wireOut_LB[53]), .outData_54(wireOut_LB[54]), .outData_55(wireOut_LB[55]), .outData_56(wireOut_LB[56]), .outData_57(wireOut_LB[57]), .outData_58(wireOut_LB[58]), .outData_59(wireOut_LB[59]), .outData_60(wireOut_LB[60]), .outData_61(wireOut_LB[61]), .outData_62(wireOut_LB[62]), .outData_63(wireOut_LB[63]), .outData_64(wireOut_LB[64]), .outData_65(wireOut_LB[65]), .outData_66(wireOut_LB[66]), .outData_67(wireOut_LB[67]), .outData_68(wireOut_LB[68]), .outData_69(wireOut_LB[69]), .outData_70(wireOut_LB[70]), .outData_71(wireOut_LB[71]), .outData_72(wireOut_LB[72]), .outData_73(wireOut_LB[73]), .outData_74(wireOut_LB[74]), .outData_75(wireOut_LB[75]), .outData_76(wireOut_LB[76]), .outData_77(wireOut_LB[77]), .outData_78(wireOut_LB[78]), .outData_79(wireOut_LB[79]), .outData_80(wireOut_LB[80]), .outData_81(wireOut_LB[81]), .outData_82(wireOut_LB[82]), .outData_83(wireOut_LB[83]), .outData_84(wireOut_LB[84]), .outData_85(wireOut_LB[85]), .outData_86(wireOut_LB[86]), .outData_87(wireOut_LB[87]), .outData_88(wireOut_LB[88]), .outData_89(wireOut_LB[89]), .outData_90(wireOut_LB[90]), .outData_91(wireOut_LB[91]), .outData_92(wireOut_LB[92]), .outData_93(wireOut_LB[93]), .outData_94(wireOut_LB[94]), .outData_95(wireOut_LB[95]), .outData_96(wireOut_LB[96]), .outData_97(wireOut_LB[97]), .outData_98(wireOut_LB[98]), .outData_99(wireOut_LB[99]), .outData_100(wireOut_LB[100]), .outData_101(wireOut_LB[101]), .outData_102(wireOut_LB[102]), .outData_103(wireOut_LB[103]), .outData_104(wireOut_LB[104]), .outData_105(wireOut_LB[105]), .outData_106(wireOut_LB[106]), .outData_107(wireOut_LB[107]), .outData_108(wireOut_LB[108]), .outData_109(wireOut_LB[109]), .outData_110(wireOut_LB[110]), .outData_111(wireOut_LB[111]), .outData_112(wireOut_LB[112]), .outData_113(wireOut_LB[113]), .outData_114(wireOut_LB[114]), .outData_115(wireOut_LB[115]), .outData_116(wireOut_LB[116]), .outData_117(wireOut_LB[117]), .outData_118(wireOut_LB[118]), .outData_119(wireOut_LB[119]), .outData_120(wireOut_LB[120]), .outData_121(wireOut_LB[121]), .outData_122(wireOut_LB[122]), .outData_123(wireOut_LB[123]), .outData_124(wireOut_LB[124]), .outData_125(wireOut_LB[125]), .outData_126(wireOut_LB[126]), .outData_127(wireOut_LB[127]), .outData_128(wireOut_LB[128]), .outData_129(wireOut_LB[129]), .outData_130(wireOut_LB[130]), .outData_131(wireOut_LB[131]), .outData_132(wireOut_LB[132]), .outData_133(wireOut_LB[133]), .outData_134(wireOut_LB[134]), .outData_135(wireOut_LB[135]), .outData_136(wireOut_LB[136]), .outData_137(wireOut_LB[137]), .outData_138(wireOut_LB[138]), .outData_139(wireOut_LB[139]), .outData_140(wireOut_LB[140]), .outData_141(wireOut_LB[141]), .outData_142(wireOut_LB[142]), .outData_143(wireOut_LB[143]), .outData_144(wireOut_LB[144]), .outData_145(wireOut_LB[145]), .outData_146(wireOut_LB[146]), .outData_147(wireOut_LB[147]), .outData_148(wireOut_LB[148]), .outData_149(wireOut_LB[149]), .outData_150(wireOut_LB[150]), .outData_151(wireOut_LB[151]), .outData_152(wireOut_LB[152]), .outData_153(wireOut_LB[153]), .outData_154(wireOut_LB[154]), .outData_155(wireOut_LB[155]), .outData_156(wireOut_LB[156]), .outData_157(wireOut_LB[157]), .outData_158(wireOut_LB[158]), .outData_159(wireOut_LB[159]), .outData_160(wireOut_LB[160]), .outData_161(wireOut_LB[161]), .outData_162(wireOut_LB[162]), .outData_163(wireOut_LB[163]), .outData_164(wireOut_LB[164]), .outData_165(wireOut_LB[165]), .outData_166(wireOut_LB[166]), .outData_167(wireOut_LB[167]), .outData_168(wireOut_LB[168]), .outData_169(wireOut_LB[169]), .outData_170(wireOut_LB[170]), .outData_171(wireOut_LB[171]), .outData_172(wireOut_LB[172]), .outData_173(wireOut_LB[173]), .outData_174(wireOut_LB[174]), .outData_175(wireOut_LB[175]), .outData_176(wireOut_LB[176]), .outData_177(wireOut_LB[177]), .outData_178(wireOut_LB[178]), .outData_179(wireOut_LB[179]), .outData_180(wireOut_LB[180]), .outData_181(wireOut_LB[181]), .outData_182(wireOut_LB[182]), .outData_183(wireOut_LB[183]), .outData_184(wireOut_LB[184]), .outData_185(wireOut_LB[185]), .outData_186(wireOut_LB[186]), .outData_187(wireOut_LB[187]), .outData_188(wireOut_LB[188]), .outData_189(wireOut_LB[189]), .outData_190(wireOut_LB[190]), .outData_191(wireOut_LB[191]), .outData_192(wireOut_LB[192]), .outData_193(wireOut_LB[193]), .outData_194(wireOut_LB[194]), .outData_195(wireOut_LB[195]), .outData_196(wireOut_LB[196]), .outData_197(wireOut_LB[197]), .outData_198(wireOut_LB[198]), .outData_199(wireOut_LB[199]), .outData_200(wireOut_LB[200]), .outData_201(wireOut_LB[201]), .outData_202(wireOut_LB[202]), .outData_203(wireOut_LB[203]), .outData_204(wireOut_LB[204]), .outData_205(wireOut_LB[205]), .outData_206(wireOut_LB[206]), .outData_207(wireOut_LB[207]), .outData_208(wireOut_LB[208]), .outData_209(wireOut_LB[209]), .outData_210(wireOut_LB[210]), .outData_211(wireOut_LB[211]), .outData_212(wireOut_LB[212]), .outData_213(wireOut_LB[213]), .outData_214(wireOut_LB[214]), .outData_215(wireOut_LB[215]), .outData_216(wireOut_LB[216]), .outData_217(wireOut_LB[217]), .outData_218(wireOut_LB[218]), .outData_219(wireOut_LB[219]), .outData_220(wireOut_LB[220]), .outData_221(wireOut_LB[221]), .outData_222(wireOut_LB[222]), .outData_223(wireOut_LB[223]), .outData_224(wireOut_LB[224]), .outData_225(wireOut_LB[225]), .outData_226(wireOut_LB[226]), .outData_227(wireOut_LB[227]), .outData_228(wireOut_LB[228]), .outData_229(wireOut_LB[229]), .outData_230(wireOut_LB[230]), .outData_231(wireOut_LB[231]), .outData_232(wireOut_LB[232]), .outData_233(wireOut_LB[233]), .outData_234(wireOut_LB[234]), .outData_235(wireOut_LB[235]), .outData_236(wireOut_LB[236]), .outData_237(wireOut_LB[237]), .outData_238(wireOut_LB[238]), .outData_239(wireOut_LB[239]), .outData_240(wireOut_LB[240]), .outData_241(wireOut_LB[241]), .outData_242(wireOut_LB[242]), .outData_243(wireOut_LB[243]), .outData_244(wireOut_LB[244]), .outData_245(wireOut_LB[245]), .outData_246(wireOut_LB[246]), .outData_247(wireOut_LB[247]), .outData_248(wireOut_LB[248]), .outData_249(wireOut_LB[249]), .outData_250(wireOut_LB[250]), .outData_251(wireOut_LB[251]), .outData_252(wireOut_LB[252]), .outData_253(wireOut_LB[253]), .outData_254(wireOut_LB[254]), .outData_255(wireOut_LB[255]), .in_start(in_start), .out_start(out_start_LB), .counter_in(counter_out_w), .clk(clk), .rst(rst));
  
  mem_stage_dp256_r mem_stage_dp256_r_inst(.inData_0(wireOut_LB[0]), .inData_1(wireOut_LB[1]), .inData_2(wireOut_LB[2]), .inData_3(wireOut_LB[3]), .inData_4(wireOut_LB[4]), .inData_5(wireOut_LB[5]), .inData_6(wireOut_LB[6]), .inData_7(wireOut_LB[7]), .inData_8(wireOut_LB[8]), .inData_9(wireOut_LB[9]), .inData_10(wireOut_LB[10]), .inData_11(wireOut_LB[11]), .inData_12(wireOut_LB[12]), .inData_13(wireOut_LB[13]), .inData_14(wireOut_LB[14]), .inData_15(wireOut_LB[15]), .inData_16(wireOut_LB[16]), .inData_17(wireOut_LB[17]), .inData_18(wireOut_LB[18]), .inData_19(wireOut_LB[19]), .inData_20(wireOut_LB[20]), .inData_21(wireOut_LB[21]), .inData_22(wireOut_LB[22]), .inData_23(wireOut_LB[23]), .inData_24(wireOut_LB[24]), .inData_25(wireOut_LB[25]), .inData_26(wireOut_LB[26]), .inData_27(wireOut_LB[27]), .inData_28(wireOut_LB[28]), .inData_29(wireOut_LB[29]), .inData_30(wireOut_LB[30]), .inData_31(wireOut_LB[31]), .inData_32(wireOut_LB[32]), .inData_33(wireOut_LB[33]), .inData_34(wireOut_LB[34]), .inData_35(wireOut_LB[35]), .inData_36(wireOut_LB[36]), .inData_37(wireOut_LB[37]), .inData_38(wireOut_LB[38]), .inData_39(wireOut_LB[39]), .inData_40(wireOut_LB[40]), .inData_41(wireOut_LB[41]), .inData_42(wireOut_LB[42]), .inData_43(wireOut_LB[43]), .inData_44(wireOut_LB[44]), .inData_45(wireOut_LB[45]), .inData_46(wireOut_LB[46]), .inData_47(wireOut_LB[47]), .inData_48(wireOut_LB[48]), .inData_49(wireOut_LB[49]), .inData_50(wireOut_LB[50]), .inData_51(wireOut_LB[51]), .inData_52(wireOut_LB[52]), .inData_53(wireOut_LB[53]), .inData_54(wireOut_LB[54]), .inData_55(wireOut_LB[55]), .inData_56(wireOut_LB[56]), .inData_57(wireOut_LB[57]), .inData_58(wireOut_LB[58]), .inData_59(wireOut_LB[59]), .inData_60(wireOut_LB[60]), .inData_61(wireOut_LB[61]), .inData_62(wireOut_LB[62]), .inData_63(wireOut_LB[63]), .inData_64(wireOut_LB[64]), .inData_65(wireOut_LB[65]), .inData_66(wireOut_LB[66]), .inData_67(wireOut_LB[67]), .inData_68(wireOut_LB[68]), .inData_69(wireOut_LB[69]), .inData_70(wireOut_LB[70]), .inData_71(wireOut_LB[71]), .inData_72(wireOut_LB[72]), .inData_73(wireOut_LB[73]), .inData_74(wireOut_LB[74]), .inData_75(wireOut_LB[75]), .inData_76(wireOut_LB[76]), .inData_77(wireOut_LB[77]), .inData_78(wireOut_LB[78]), .inData_79(wireOut_LB[79]), .inData_80(wireOut_LB[80]), .inData_81(wireOut_LB[81]), .inData_82(wireOut_LB[82]), .inData_83(wireOut_LB[83]), .inData_84(wireOut_LB[84]), .inData_85(wireOut_LB[85]), .inData_86(wireOut_LB[86]), .inData_87(wireOut_LB[87]), .inData_88(wireOut_LB[88]), .inData_89(wireOut_LB[89]), .inData_90(wireOut_LB[90]), .inData_91(wireOut_LB[91]), .inData_92(wireOut_LB[92]), .inData_93(wireOut_LB[93]), .inData_94(wireOut_LB[94]), .inData_95(wireOut_LB[95]), .inData_96(wireOut_LB[96]), .inData_97(wireOut_LB[97]), .inData_98(wireOut_LB[98]), .inData_99(wireOut_LB[99]), .inData_100(wireOut_LB[100]), .inData_101(wireOut_LB[101]), .inData_102(wireOut_LB[102]), .inData_103(wireOut_LB[103]), .inData_104(wireOut_LB[104]), .inData_105(wireOut_LB[105]), .inData_106(wireOut_LB[106]), .inData_107(wireOut_LB[107]), .inData_108(wireOut_LB[108]), .inData_109(wireOut_LB[109]), .inData_110(wireOut_LB[110]), .inData_111(wireOut_LB[111]), .inData_112(wireOut_LB[112]), .inData_113(wireOut_LB[113]), .inData_114(wireOut_LB[114]), .inData_115(wireOut_LB[115]), .inData_116(wireOut_LB[116]), .inData_117(wireOut_LB[117]), .inData_118(wireOut_LB[118]), .inData_119(wireOut_LB[119]), .inData_120(wireOut_LB[120]), .inData_121(wireOut_LB[121]), .inData_122(wireOut_LB[122]), .inData_123(wireOut_LB[123]), .inData_124(wireOut_LB[124]), .inData_125(wireOut_LB[125]), .inData_126(wireOut_LB[126]), .inData_127(wireOut_LB[127]), .inData_128(wireOut_LB[128]), .inData_129(wireOut_LB[129]), .inData_130(wireOut_LB[130]), .inData_131(wireOut_LB[131]), .inData_132(wireOut_LB[132]), .inData_133(wireOut_LB[133]), .inData_134(wireOut_LB[134]), .inData_135(wireOut_LB[135]), .inData_136(wireOut_LB[136]), .inData_137(wireOut_LB[137]), .inData_138(wireOut_LB[138]), .inData_139(wireOut_LB[139]), .inData_140(wireOut_LB[140]), .inData_141(wireOut_LB[141]), .inData_142(wireOut_LB[142]), .inData_143(wireOut_LB[143]), .inData_144(wireOut_LB[144]), .inData_145(wireOut_LB[145]), .inData_146(wireOut_LB[146]), .inData_147(wireOut_LB[147]), .inData_148(wireOut_LB[148]), .inData_149(wireOut_LB[149]), .inData_150(wireOut_LB[150]), .inData_151(wireOut_LB[151]), .inData_152(wireOut_LB[152]), .inData_153(wireOut_LB[153]), .inData_154(wireOut_LB[154]), .inData_155(wireOut_LB[155]), .inData_156(wireOut_LB[156]), .inData_157(wireOut_LB[157]), .inData_158(wireOut_LB[158]), .inData_159(wireOut_LB[159]), .inData_160(wireOut_LB[160]), .inData_161(wireOut_LB[161]), .inData_162(wireOut_LB[162]), .inData_163(wireOut_LB[163]), .inData_164(wireOut_LB[164]), .inData_165(wireOut_LB[165]), .inData_166(wireOut_LB[166]), .inData_167(wireOut_LB[167]), .inData_168(wireOut_LB[168]), .inData_169(wireOut_LB[169]), .inData_170(wireOut_LB[170]), .inData_171(wireOut_LB[171]), .inData_172(wireOut_LB[172]), .inData_173(wireOut_LB[173]), .inData_174(wireOut_LB[174]), .inData_175(wireOut_LB[175]), .inData_176(wireOut_LB[176]), .inData_177(wireOut_LB[177]), .inData_178(wireOut_LB[178]), .inData_179(wireOut_LB[179]), .inData_180(wireOut_LB[180]), .inData_181(wireOut_LB[181]), .inData_182(wireOut_LB[182]), .inData_183(wireOut_LB[183]), .inData_184(wireOut_LB[184]), .inData_185(wireOut_LB[185]), .inData_186(wireOut_LB[186]), .inData_187(wireOut_LB[187]), .inData_188(wireOut_LB[188]), .inData_189(wireOut_LB[189]), .inData_190(wireOut_LB[190]), .inData_191(wireOut_LB[191]), .inData_192(wireOut_LB[192]), .inData_193(wireOut_LB[193]), .inData_194(wireOut_LB[194]), .inData_195(wireOut_LB[195]), .inData_196(wireOut_LB[196]), .inData_197(wireOut_LB[197]), .inData_198(wireOut_LB[198]), .inData_199(wireOut_LB[199]), .inData_200(wireOut_LB[200]), .inData_201(wireOut_LB[201]), .inData_202(wireOut_LB[202]), .inData_203(wireOut_LB[203]), .inData_204(wireOut_LB[204]), .inData_205(wireOut_LB[205]), .inData_206(wireOut_LB[206]), .inData_207(wireOut_LB[207]), .inData_208(wireOut_LB[208]), .inData_209(wireOut_LB[209]), .inData_210(wireOut_LB[210]), .inData_211(wireOut_LB[211]), .inData_212(wireOut_LB[212]), .inData_213(wireOut_LB[213]), .inData_214(wireOut_LB[214]), .inData_215(wireOut_LB[215]), .inData_216(wireOut_LB[216]), .inData_217(wireOut_LB[217]), .inData_218(wireOut_LB[218]), .inData_219(wireOut_LB[219]), .inData_220(wireOut_LB[220]), .inData_221(wireOut_LB[221]), .inData_222(wireOut_LB[222]), .inData_223(wireOut_LB[223]), .inData_224(wireOut_LB[224]), .inData_225(wireOut_LB[225]), .inData_226(wireOut_LB[226]), .inData_227(wireOut_LB[227]), .inData_228(wireOut_LB[228]), .inData_229(wireOut_LB[229]), .inData_230(wireOut_LB[230]), .inData_231(wireOut_LB[231]), .inData_232(wireOut_LB[232]), .inData_233(wireOut_LB[233]), .inData_234(wireOut_LB[234]), .inData_235(wireOut_LB[235]), .inData_236(wireOut_LB[236]), .inData_237(wireOut_LB[237]), .inData_238(wireOut_LB[238]), .inData_239(wireOut_LB[239]), .inData_240(wireOut_LB[240]), .inData_241(wireOut_LB[241]), .inData_242(wireOut_LB[242]), .inData_243(wireOut_LB[243]), .inData_244(wireOut_LB[244]), .inData_245(wireOut_LB[245]), .inData_246(wireOut_LB[246]), .inData_247(wireOut_LB[247]), .inData_248(wireOut_LB[248]), .inData_249(wireOut_LB[249]), .inData_250(wireOut_LB[250]), .inData_251(wireOut_LB[251]), .inData_252(wireOut_LB[252]), .inData_253(wireOut_LB[253]), .inData_254(wireOut_LB[254]), .inData_255(wireOut_LB[255]), .outData_0(wireIn_RB[0]), .outData_1(wireIn_RB[1]), .outData_2(wireIn_RB[2]), .outData_3(wireIn_RB[3]), .outData_4(wireIn_RB[4]), .outData_5(wireIn_RB[5]), .outData_6(wireIn_RB[6]), .outData_7(wireIn_RB[7]), .outData_8(wireIn_RB[8]), .outData_9(wireIn_RB[9]), .outData_10(wireIn_RB[10]), .outData_11(wireIn_RB[11]), .outData_12(wireIn_RB[12]), .outData_13(wireIn_RB[13]), .outData_14(wireIn_RB[14]), .outData_15(wireIn_RB[15]), .outData_16(wireIn_RB[16]), .outData_17(wireIn_RB[17]), .outData_18(wireIn_RB[18]), .outData_19(wireIn_RB[19]), .outData_20(wireIn_RB[20]), .outData_21(wireIn_RB[21]), .outData_22(wireIn_RB[22]), .outData_23(wireIn_RB[23]), .outData_24(wireIn_RB[24]), .outData_25(wireIn_RB[25]), .outData_26(wireIn_RB[26]), .outData_27(wireIn_RB[27]), .outData_28(wireIn_RB[28]), .outData_29(wireIn_RB[29]), .outData_30(wireIn_RB[30]), .outData_31(wireIn_RB[31]), .outData_32(wireIn_RB[32]), .outData_33(wireIn_RB[33]), .outData_34(wireIn_RB[34]), .outData_35(wireIn_RB[35]), .outData_36(wireIn_RB[36]), .outData_37(wireIn_RB[37]), .outData_38(wireIn_RB[38]), .outData_39(wireIn_RB[39]), .outData_40(wireIn_RB[40]), .outData_41(wireIn_RB[41]), .outData_42(wireIn_RB[42]), .outData_43(wireIn_RB[43]), .outData_44(wireIn_RB[44]), .outData_45(wireIn_RB[45]), .outData_46(wireIn_RB[46]), .outData_47(wireIn_RB[47]), .outData_48(wireIn_RB[48]), .outData_49(wireIn_RB[49]), .outData_50(wireIn_RB[50]), .outData_51(wireIn_RB[51]), .outData_52(wireIn_RB[52]), .outData_53(wireIn_RB[53]), .outData_54(wireIn_RB[54]), .outData_55(wireIn_RB[55]), .outData_56(wireIn_RB[56]), .outData_57(wireIn_RB[57]), .outData_58(wireIn_RB[58]), .outData_59(wireIn_RB[59]), .outData_60(wireIn_RB[60]), .outData_61(wireIn_RB[61]), .outData_62(wireIn_RB[62]), .outData_63(wireIn_RB[63]), .outData_64(wireIn_RB[64]), .outData_65(wireIn_RB[65]), .outData_66(wireIn_RB[66]), .outData_67(wireIn_RB[67]), .outData_68(wireIn_RB[68]), .outData_69(wireIn_RB[69]), .outData_70(wireIn_RB[70]), .outData_71(wireIn_RB[71]), .outData_72(wireIn_RB[72]), .outData_73(wireIn_RB[73]), .outData_74(wireIn_RB[74]), .outData_75(wireIn_RB[75]), .outData_76(wireIn_RB[76]), .outData_77(wireIn_RB[77]), .outData_78(wireIn_RB[78]), .outData_79(wireIn_RB[79]), .outData_80(wireIn_RB[80]), .outData_81(wireIn_RB[81]), .outData_82(wireIn_RB[82]), .outData_83(wireIn_RB[83]), .outData_84(wireIn_RB[84]), .outData_85(wireIn_RB[85]), .outData_86(wireIn_RB[86]), .outData_87(wireIn_RB[87]), .outData_88(wireIn_RB[88]), .outData_89(wireIn_RB[89]), .outData_90(wireIn_RB[90]), .outData_91(wireIn_RB[91]), .outData_92(wireIn_RB[92]), .outData_93(wireIn_RB[93]), .outData_94(wireIn_RB[94]), .outData_95(wireIn_RB[95]), .outData_96(wireIn_RB[96]), .outData_97(wireIn_RB[97]), .outData_98(wireIn_RB[98]), .outData_99(wireIn_RB[99]), .outData_100(wireIn_RB[100]), .outData_101(wireIn_RB[101]), .outData_102(wireIn_RB[102]), .outData_103(wireIn_RB[103]), .outData_104(wireIn_RB[104]), .outData_105(wireIn_RB[105]), .outData_106(wireIn_RB[106]), .outData_107(wireIn_RB[107]), .outData_108(wireIn_RB[108]), .outData_109(wireIn_RB[109]), .outData_110(wireIn_RB[110]), .outData_111(wireIn_RB[111]), .outData_112(wireIn_RB[112]), .outData_113(wireIn_RB[113]), .outData_114(wireIn_RB[114]), .outData_115(wireIn_RB[115]), .outData_116(wireIn_RB[116]), .outData_117(wireIn_RB[117]), .outData_118(wireIn_RB[118]), .outData_119(wireIn_RB[119]), .outData_120(wireIn_RB[120]), .outData_121(wireIn_RB[121]), .outData_122(wireIn_RB[122]), .outData_123(wireIn_RB[123]), .outData_124(wireIn_RB[124]), .outData_125(wireIn_RB[125]), .outData_126(wireIn_RB[126]), .outData_127(wireIn_RB[127]), .outData_128(wireIn_RB[128]), .outData_129(wireIn_RB[129]), .outData_130(wireIn_RB[130]), .outData_131(wireIn_RB[131]), .outData_132(wireIn_RB[132]), .outData_133(wireIn_RB[133]), .outData_134(wireIn_RB[134]), .outData_135(wireIn_RB[135]), .outData_136(wireIn_RB[136]), .outData_137(wireIn_RB[137]), .outData_138(wireIn_RB[138]), .outData_139(wireIn_RB[139]), .outData_140(wireIn_RB[140]), .outData_141(wireIn_RB[141]), .outData_142(wireIn_RB[142]), .outData_143(wireIn_RB[143]), .outData_144(wireIn_RB[144]), .outData_145(wireIn_RB[145]), .outData_146(wireIn_RB[146]), .outData_147(wireIn_RB[147]), .outData_148(wireIn_RB[148]), .outData_149(wireIn_RB[149]), .outData_150(wireIn_RB[150]), .outData_151(wireIn_RB[151]), .outData_152(wireIn_RB[152]), .outData_153(wireIn_RB[153]), .outData_154(wireIn_RB[154]), .outData_155(wireIn_RB[155]), .outData_156(wireIn_RB[156]), .outData_157(wireIn_RB[157]), .outData_158(wireIn_RB[158]), .outData_159(wireIn_RB[159]), .outData_160(wireIn_RB[160]), .outData_161(wireIn_RB[161]), .outData_162(wireIn_RB[162]), .outData_163(wireIn_RB[163]), .outData_164(wireIn_RB[164]), .outData_165(wireIn_RB[165]), .outData_166(wireIn_RB[166]), .outData_167(wireIn_RB[167]), .outData_168(wireIn_RB[168]), .outData_169(wireIn_RB[169]), .outData_170(wireIn_RB[170]), .outData_171(wireIn_RB[171]), .outData_172(wireIn_RB[172]), .outData_173(wireIn_RB[173]), .outData_174(wireIn_RB[174]), .outData_175(wireIn_RB[175]), .outData_176(wireIn_RB[176]), .outData_177(wireIn_RB[177]), .outData_178(wireIn_RB[178]), .outData_179(wireIn_RB[179]), .outData_180(wireIn_RB[180]), .outData_181(wireIn_RB[181]), .outData_182(wireIn_RB[182]), .outData_183(wireIn_RB[183]), .outData_184(wireIn_RB[184]), .outData_185(wireIn_RB[185]), .outData_186(wireIn_RB[186]), .outData_187(wireIn_RB[187]), .outData_188(wireIn_RB[188]), .outData_189(wireIn_RB[189]), .outData_190(wireIn_RB[190]), .outData_191(wireIn_RB[191]), .outData_192(wireIn_RB[192]), .outData_193(wireIn_RB[193]), .outData_194(wireIn_RB[194]), .outData_195(wireIn_RB[195]), .outData_196(wireIn_RB[196]), .outData_197(wireIn_RB[197]), .outData_198(wireIn_RB[198]), .outData_199(wireIn_RB[199]), .outData_200(wireIn_RB[200]), .outData_201(wireIn_RB[201]), .outData_202(wireIn_RB[202]), .outData_203(wireIn_RB[203]), .outData_204(wireIn_RB[204]), .outData_205(wireIn_RB[205]), .outData_206(wireIn_RB[206]), .outData_207(wireIn_RB[207]), .outData_208(wireIn_RB[208]), .outData_209(wireIn_RB[209]), .outData_210(wireIn_RB[210]), .outData_211(wireIn_RB[211]), .outData_212(wireIn_RB[212]), .outData_213(wireIn_RB[213]), .outData_214(wireIn_RB[214]), .outData_215(wireIn_RB[215]), .outData_216(wireIn_RB[216]), .outData_217(wireIn_RB[217]), .outData_218(wireIn_RB[218]), .outData_219(wireIn_RB[219]), .outData_220(wireIn_RB[220]), .outData_221(wireIn_RB[221]), .outData_222(wireIn_RB[222]), .outData_223(wireIn_RB[223]), .outData_224(wireIn_RB[224]), .outData_225(wireIn_RB[225]), .outData_226(wireIn_RB[226]), .outData_227(wireIn_RB[227]), .outData_228(wireIn_RB[228]), .outData_229(wireIn_RB[229]), .outData_230(wireIn_RB[230]), .outData_231(wireIn_RB[231]), .outData_232(wireIn_RB[232]), .outData_233(wireIn_RB[233]), .outData_234(wireIn_RB[234]), .outData_235(wireIn_RB[235]), .outData_236(wireIn_RB[236]), .outData_237(wireIn_RB[237]), .outData_238(wireIn_RB[238]), .outData_239(wireIn_RB[239]), .outData_240(wireIn_RB[240]), .outData_241(wireIn_RB[241]), .outData_242(wireIn_RB[242]), .outData_243(wireIn_RB[243]), .outData_244(wireIn_RB[244]), .outData_245(wireIn_RB[245]), .outData_246(wireIn_RB[246]), .outData_247(wireIn_RB[247]), .outData_248(wireIn_RB[248]), .outData_249(wireIn_RB[249]), .outData_250(wireIn_RB[250]), .outData_251(wireIn_RB[251]), .outData_252(wireIn_RB[252]), .outData_253(wireIn_RB[253]), .outData_254(wireIn_RB[254]), .outData_255(wireIn_RB[255]), .in_start(out_start_LB), .out_start(out_start_MemStage), .clk(clk), 
 .counter_in(counter_out_w), .rst(rst));
  
  egressStage_p256 egressStage_p256_inst(.inData_0(wireIn_RB[0]), .inData_1(wireIn_RB[1]), .inData_2(wireIn_RB[2]), .inData_3(wireIn_RB[3]), .inData_4(wireIn_RB[4]), .inData_5(wireIn_RB[5]), .inData_6(wireIn_RB[6]), .inData_7(wireIn_RB[7]), .inData_8(wireIn_RB[8]), .inData_9(wireIn_RB[9]), .inData_10(wireIn_RB[10]), .inData_11(wireIn_RB[11]), .inData_12(wireIn_RB[12]), .inData_13(wireIn_RB[13]), .inData_14(wireIn_RB[14]), .inData_15(wireIn_RB[15]), .inData_16(wireIn_RB[16]), .inData_17(wireIn_RB[17]), .inData_18(wireIn_RB[18]), .inData_19(wireIn_RB[19]), .inData_20(wireIn_RB[20]), .inData_21(wireIn_RB[21]), .inData_22(wireIn_RB[22]), .inData_23(wireIn_RB[23]), .inData_24(wireIn_RB[24]), .inData_25(wireIn_RB[25]), .inData_26(wireIn_RB[26]), .inData_27(wireIn_RB[27]), .inData_28(wireIn_RB[28]), .inData_29(wireIn_RB[29]), .inData_30(wireIn_RB[30]), .inData_31(wireIn_RB[31]), .inData_32(wireIn_RB[32]), .inData_33(wireIn_RB[33]), .inData_34(wireIn_RB[34]), .inData_35(wireIn_RB[35]), .inData_36(wireIn_RB[36]), .inData_37(wireIn_RB[37]), .inData_38(wireIn_RB[38]), .inData_39(wireIn_RB[39]), .inData_40(wireIn_RB[40]), .inData_41(wireIn_RB[41]), .inData_42(wireIn_RB[42]), .inData_43(wireIn_RB[43]), .inData_44(wireIn_RB[44]), .inData_45(wireIn_RB[45]), .inData_46(wireIn_RB[46]), .inData_47(wireIn_RB[47]), .inData_48(wireIn_RB[48]), .inData_49(wireIn_RB[49]), .inData_50(wireIn_RB[50]), .inData_51(wireIn_RB[51]), .inData_52(wireIn_RB[52]), .inData_53(wireIn_RB[53]), .inData_54(wireIn_RB[54]), .inData_55(wireIn_RB[55]), .inData_56(wireIn_RB[56]), .inData_57(wireIn_RB[57]), .inData_58(wireIn_RB[58]), .inData_59(wireIn_RB[59]), .inData_60(wireIn_RB[60]), .inData_61(wireIn_RB[61]), .inData_62(wireIn_RB[62]), .inData_63(wireIn_RB[63]), .inData_64(wireIn_RB[64]), .inData_65(wireIn_RB[65]), .inData_66(wireIn_RB[66]), .inData_67(wireIn_RB[67]), .inData_68(wireIn_RB[68]), .inData_69(wireIn_RB[69]), .inData_70(wireIn_RB[70]), .inData_71(wireIn_RB[71]), .inData_72(wireIn_RB[72]), .inData_73(wireIn_RB[73]), .inData_74(wireIn_RB[74]), .inData_75(wireIn_RB[75]), .inData_76(wireIn_RB[76]), .inData_77(wireIn_RB[77]), .inData_78(wireIn_RB[78]), .inData_79(wireIn_RB[79]), .inData_80(wireIn_RB[80]), .inData_81(wireIn_RB[81]), .inData_82(wireIn_RB[82]), .inData_83(wireIn_RB[83]), .inData_84(wireIn_RB[84]), .inData_85(wireIn_RB[85]), .inData_86(wireIn_RB[86]), .inData_87(wireIn_RB[87]), .inData_88(wireIn_RB[88]), .inData_89(wireIn_RB[89]), .inData_90(wireIn_RB[90]), .inData_91(wireIn_RB[91]), .inData_92(wireIn_RB[92]), .inData_93(wireIn_RB[93]), .inData_94(wireIn_RB[94]), .inData_95(wireIn_RB[95]), .inData_96(wireIn_RB[96]), .inData_97(wireIn_RB[97]), .inData_98(wireIn_RB[98]), .inData_99(wireIn_RB[99]), .inData_100(wireIn_RB[100]), .inData_101(wireIn_RB[101]), .inData_102(wireIn_RB[102]), .inData_103(wireIn_RB[103]), .inData_104(wireIn_RB[104]), .inData_105(wireIn_RB[105]), .inData_106(wireIn_RB[106]), .inData_107(wireIn_RB[107]), .inData_108(wireIn_RB[108]), .inData_109(wireIn_RB[109]), .inData_110(wireIn_RB[110]), .inData_111(wireIn_RB[111]), .inData_112(wireIn_RB[112]), .inData_113(wireIn_RB[113]), .inData_114(wireIn_RB[114]), .inData_115(wireIn_RB[115]), .inData_116(wireIn_RB[116]), .inData_117(wireIn_RB[117]), .inData_118(wireIn_RB[118]), .inData_119(wireIn_RB[119]), .inData_120(wireIn_RB[120]), .inData_121(wireIn_RB[121]), .inData_122(wireIn_RB[122]), .inData_123(wireIn_RB[123]), .inData_124(wireIn_RB[124]), .inData_125(wireIn_RB[125]), .inData_126(wireIn_RB[126]), .inData_127(wireIn_RB[127]), .inData_128(wireIn_RB[128]), .inData_129(wireIn_RB[129]), .inData_130(wireIn_RB[130]), .inData_131(wireIn_RB[131]), .inData_132(wireIn_RB[132]), .inData_133(wireIn_RB[133]), .inData_134(wireIn_RB[134]), .inData_135(wireIn_RB[135]), .inData_136(wireIn_RB[136]), .inData_137(wireIn_RB[137]), .inData_138(wireIn_RB[138]), .inData_139(wireIn_RB[139]), .inData_140(wireIn_RB[140]), .inData_141(wireIn_RB[141]), .inData_142(wireIn_RB[142]), .inData_143(wireIn_RB[143]), .inData_144(wireIn_RB[144]), .inData_145(wireIn_RB[145]), .inData_146(wireIn_RB[146]), .inData_147(wireIn_RB[147]), .inData_148(wireIn_RB[148]), .inData_149(wireIn_RB[149]), .inData_150(wireIn_RB[150]), .inData_151(wireIn_RB[151]), .inData_152(wireIn_RB[152]), .inData_153(wireIn_RB[153]), .inData_154(wireIn_RB[154]), .inData_155(wireIn_RB[155]), .inData_156(wireIn_RB[156]), .inData_157(wireIn_RB[157]), .inData_158(wireIn_RB[158]), .inData_159(wireIn_RB[159]), .inData_160(wireIn_RB[160]), .inData_161(wireIn_RB[161]), .inData_162(wireIn_RB[162]), .inData_163(wireIn_RB[163]), .inData_164(wireIn_RB[164]), .inData_165(wireIn_RB[165]), .inData_166(wireIn_RB[166]), .inData_167(wireIn_RB[167]), .inData_168(wireIn_RB[168]), .inData_169(wireIn_RB[169]), .inData_170(wireIn_RB[170]), .inData_171(wireIn_RB[171]), .inData_172(wireIn_RB[172]), .inData_173(wireIn_RB[173]), .inData_174(wireIn_RB[174]), .inData_175(wireIn_RB[175]), .inData_176(wireIn_RB[176]), .inData_177(wireIn_RB[177]), .inData_178(wireIn_RB[178]), .inData_179(wireIn_RB[179]), .inData_180(wireIn_RB[180]), .inData_181(wireIn_RB[181]), .inData_182(wireIn_RB[182]), .inData_183(wireIn_RB[183]), .inData_184(wireIn_RB[184]), .inData_185(wireIn_RB[185]), .inData_186(wireIn_RB[186]), .inData_187(wireIn_RB[187]), .inData_188(wireIn_RB[188]), .inData_189(wireIn_RB[189]), .inData_190(wireIn_RB[190]), .inData_191(wireIn_RB[191]), .inData_192(wireIn_RB[192]), .inData_193(wireIn_RB[193]), .inData_194(wireIn_RB[194]), .inData_195(wireIn_RB[195]), .inData_196(wireIn_RB[196]), .inData_197(wireIn_RB[197]), .inData_198(wireIn_RB[198]), .inData_199(wireIn_RB[199]), .inData_200(wireIn_RB[200]), .inData_201(wireIn_RB[201]), .inData_202(wireIn_RB[202]), .inData_203(wireIn_RB[203]), .inData_204(wireIn_RB[204]), .inData_205(wireIn_RB[205]), .inData_206(wireIn_RB[206]), .inData_207(wireIn_RB[207]), .inData_208(wireIn_RB[208]), .inData_209(wireIn_RB[209]), .inData_210(wireIn_RB[210]), .inData_211(wireIn_RB[211]), .inData_212(wireIn_RB[212]), .inData_213(wireIn_RB[213]), .inData_214(wireIn_RB[214]), .inData_215(wireIn_RB[215]), .inData_216(wireIn_RB[216]), .inData_217(wireIn_RB[217]), .inData_218(wireIn_RB[218]), .inData_219(wireIn_RB[219]), .inData_220(wireIn_RB[220]), .inData_221(wireIn_RB[221]), .inData_222(wireIn_RB[222]), .inData_223(wireIn_RB[223]), .inData_224(wireIn_RB[224]), .inData_225(wireIn_RB[225]), .inData_226(wireIn_RB[226]), .inData_227(wireIn_RB[227]), .inData_228(wireIn_RB[228]), .inData_229(wireIn_RB[229]), .inData_230(wireIn_RB[230]), .inData_231(wireIn_RB[231]), .inData_232(wireIn_RB[232]), .inData_233(wireIn_RB[233]), .inData_234(wireIn_RB[234]), .inData_235(wireIn_RB[235]), .inData_236(wireIn_RB[236]), .inData_237(wireIn_RB[237]), .inData_238(wireIn_RB[238]), .inData_239(wireIn_RB[239]), .inData_240(wireIn_RB[240]), .inData_241(wireIn_RB[241]), .inData_242(wireIn_RB[242]), .inData_243(wireIn_RB[243]), .inData_244(wireIn_RB[244]), .inData_245(wireIn_RB[245]), .inData_246(wireIn_RB[246]), .inData_247(wireIn_RB[247]), .inData_248(wireIn_RB[248]), .inData_249(wireIn_RB[249]), .inData_250(wireIn_RB[250]), .inData_251(wireIn_RB[251]), .inData_252(wireIn_RB[252]), .inData_253(wireIn_RB[253]), .inData_254(wireIn_RB[254]), .inData_255(wireIn_RB[255]), .outData_0(wireOut[0]), .outData_1(wireOut[1]), .outData_2(wireOut[2]), .outData_3(wireOut[3]), .outData_4(wireOut[4]), .outData_5(wireOut[5]), .outData_6(wireOut[6]), .outData_7(wireOut[7]), .outData_8(wireOut[8]), .outData_9(wireOut[9]), .outData_10(wireOut[10]), .outData_11(wireOut[11]), .outData_12(wireOut[12]), .outData_13(wireOut[13]), .outData_14(wireOut[14]), .outData_15(wireOut[15]), .outData_16(wireOut[16]), .outData_17(wireOut[17]), .outData_18(wireOut[18]), .outData_19(wireOut[19]), .outData_20(wireOut[20]), .outData_21(wireOut[21]), .outData_22(wireOut[22]), .outData_23(wireOut[23]), .outData_24(wireOut[24]), .outData_25(wireOut[25]), .outData_26(wireOut[26]), .outData_27(wireOut[27]), .outData_28(wireOut[28]), .outData_29(wireOut[29]), .outData_30(wireOut[30]), .outData_31(wireOut[31]), .outData_32(wireOut[32]), .outData_33(wireOut[33]), .outData_34(wireOut[34]), .outData_35(wireOut[35]), .outData_36(wireOut[36]), .outData_37(wireOut[37]), .outData_38(wireOut[38]), .outData_39(wireOut[39]), .outData_40(wireOut[40]), .outData_41(wireOut[41]), .outData_42(wireOut[42]), .outData_43(wireOut[43]), .outData_44(wireOut[44]), .outData_45(wireOut[45]), .outData_46(wireOut[46]), .outData_47(wireOut[47]), .outData_48(wireOut[48]), .outData_49(wireOut[49]), .outData_50(wireOut[50]), .outData_51(wireOut[51]), .outData_52(wireOut[52]), .outData_53(wireOut[53]), .outData_54(wireOut[54]), .outData_55(wireOut[55]), .outData_56(wireOut[56]), .outData_57(wireOut[57]), .outData_58(wireOut[58]), .outData_59(wireOut[59]), .outData_60(wireOut[60]), .outData_61(wireOut[61]), .outData_62(wireOut[62]), .outData_63(wireOut[63]), .outData_64(wireOut[64]), .outData_65(wireOut[65]), .outData_66(wireOut[66]), .outData_67(wireOut[67]), .outData_68(wireOut[68]), .outData_69(wireOut[69]), .outData_70(wireOut[70]), .outData_71(wireOut[71]), .outData_72(wireOut[72]), .outData_73(wireOut[73]), .outData_74(wireOut[74]), .outData_75(wireOut[75]), .outData_76(wireOut[76]), .outData_77(wireOut[77]), .outData_78(wireOut[78]), .outData_79(wireOut[79]), .outData_80(wireOut[80]), .outData_81(wireOut[81]), .outData_82(wireOut[82]), .outData_83(wireOut[83]), .outData_84(wireOut[84]), .outData_85(wireOut[85]), .outData_86(wireOut[86]), .outData_87(wireOut[87]), .outData_88(wireOut[88]), .outData_89(wireOut[89]), .outData_90(wireOut[90]), .outData_91(wireOut[91]), .outData_92(wireOut[92]), .outData_93(wireOut[93]), .outData_94(wireOut[94]), .outData_95(wireOut[95]), .outData_96(wireOut[96]), .outData_97(wireOut[97]), .outData_98(wireOut[98]), .outData_99(wireOut[99]), .outData_100(wireOut[100]), .outData_101(wireOut[101]), .outData_102(wireOut[102]), .outData_103(wireOut[103]), .outData_104(wireOut[104]), .outData_105(wireOut[105]), .outData_106(wireOut[106]), .outData_107(wireOut[107]), .outData_108(wireOut[108]), .outData_109(wireOut[109]), .outData_110(wireOut[110]), .outData_111(wireOut[111]), .outData_112(wireOut[112]), .outData_113(wireOut[113]), .outData_114(wireOut[114]), .outData_115(wireOut[115]), .outData_116(wireOut[116]), .outData_117(wireOut[117]), .outData_118(wireOut[118]), .outData_119(wireOut[119]), .outData_120(wireOut[120]), .outData_121(wireOut[121]), .outData_122(wireOut[122]), .outData_123(wireOut[123]), .outData_124(wireOut[124]), .outData_125(wireOut[125]), .outData_126(wireOut[126]), .outData_127(wireOut[127]), .outData_128(wireOut[128]), .outData_129(wireOut[129]), .outData_130(wireOut[130]), .outData_131(wireOut[131]), .outData_132(wireOut[132]), .outData_133(wireOut[133]), .outData_134(wireOut[134]), .outData_135(wireOut[135]), .outData_136(wireOut[136]), .outData_137(wireOut[137]), .outData_138(wireOut[138]), .outData_139(wireOut[139]), .outData_140(wireOut[140]), .outData_141(wireOut[141]), .outData_142(wireOut[142]), .outData_143(wireOut[143]), .outData_144(wireOut[144]), .outData_145(wireOut[145]), .outData_146(wireOut[146]), .outData_147(wireOut[147]), .outData_148(wireOut[148]), .outData_149(wireOut[149]), .outData_150(wireOut[150]), .outData_151(wireOut[151]), .outData_152(wireOut[152]), .outData_153(wireOut[153]), .outData_154(wireOut[154]), .outData_155(wireOut[155]), .outData_156(wireOut[156]), .outData_157(wireOut[157]), .outData_158(wireOut[158]), .outData_159(wireOut[159]), .outData_160(wireOut[160]), .outData_161(wireOut[161]), .outData_162(wireOut[162]), .outData_163(wireOut[163]), .outData_164(wireOut[164]), .outData_165(wireOut[165]), .outData_166(wireOut[166]), .outData_167(wireOut[167]), .outData_168(wireOut[168]), .outData_169(wireOut[169]), .outData_170(wireOut[170]), .outData_171(wireOut[171]), .outData_172(wireOut[172]), .outData_173(wireOut[173]), .outData_174(wireOut[174]), .outData_175(wireOut[175]), .outData_176(wireOut[176]), .outData_177(wireOut[177]), .outData_178(wireOut[178]), .outData_179(wireOut[179]), .outData_180(wireOut[180]), .outData_181(wireOut[181]), .outData_182(wireOut[182]), .outData_183(wireOut[183]), .outData_184(wireOut[184]), .outData_185(wireOut[185]), .outData_186(wireOut[186]), .outData_187(wireOut[187]), .outData_188(wireOut[188]), .outData_189(wireOut[189]), .outData_190(wireOut[190]), .outData_191(wireOut[191]), .outData_192(wireOut[192]), .outData_193(wireOut[193]), .outData_194(wireOut[194]), .outData_195(wireOut[195]), .outData_196(wireOut[196]), .outData_197(wireOut[197]), .outData_198(wireOut[198]), .outData_199(wireOut[199]), .outData_200(wireOut[200]), .outData_201(wireOut[201]), .outData_202(wireOut[202]), .outData_203(wireOut[203]), .outData_204(wireOut[204]), .outData_205(wireOut[205]), .outData_206(wireOut[206]), .outData_207(wireOut[207]), .outData_208(wireOut[208]), .outData_209(wireOut[209]), .outData_210(wireOut[210]), .outData_211(wireOut[211]), .outData_212(wireOut[212]), .outData_213(wireOut[213]), .outData_214(wireOut[214]), .outData_215(wireOut[215]), .outData_216(wireOut[216]), .outData_217(wireOut[217]), .outData_218(wireOut[218]), .outData_219(wireOut[219]), .outData_220(wireOut[220]), .outData_221(wireOut[221]), .outData_222(wireOut[222]), .outData_223(wireOut[223]), .outData_224(wireOut[224]), .outData_225(wireOut[225]), .outData_226(wireOut[226]), .outData_227(wireOut[227]), .outData_228(wireOut[228]), .outData_229(wireOut[229]), .outData_230(wireOut[230]), .outData_231(wireOut[231]), .outData_232(wireOut[232]), .outData_233(wireOut[233]), .outData_234(wireOut[234]), .outData_235(wireOut[235]), .outData_236(wireOut[236]), .outData_237(wireOut[237]), .outData_238(wireOut[238]), .outData_239(wireOut[239]), .outData_240(wireOut[240]), .outData_241(wireOut[241]), .outData_242(wireOut[242]), .outData_243(wireOut[243]), .outData_244(wireOut[244]), .outData_245(wireOut[245]), .outData_246(wireOut[246]), .outData_247(wireOut[247]), .outData_248(wireOut[248]), .outData_249(wireOut[249]), .outData_250(wireOut[250]), .outData_251(wireOut[251]), .outData_252(wireOut[252]), .outData_253(wireOut[253]), .outData_254(wireOut[254]), .outData_255(wireOut[255]), .in_start(out_start_MemStage), .out_start(out_start_RB), .counter_in(counter_out_w), .clk(clk), .rst(rst));
  
  
  always@(posedge clk)             
  begin                            
    if(rst) begin                    
      outData_0 <= 0;    
      outData_1 <= 0;    
      outData_2 <= 0;    
      outData_3 <= 0;    
      outData_4 <= 0;    
      outData_5 <= 0;    
      outData_6 <= 0;    
      outData_7 <= 0;    
      outData_8 <= 0;    
      outData_9 <= 0;    
      outData_10 <= 0;    
      outData_11 <= 0;    
      outData_12 <= 0;    
      outData_13 <= 0;    
      outData_14 <= 0;    
      outData_15 <= 0;    
      outData_16 <= 0;    
      outData_17 <= 0;    
      outData_18 <= 0;    
      outData_19 <= 0;    
      outData_20 <= 0;    
      outData_21 <= 0;    
      outData_22 <= 0;    
      outData_23 <= 0;    
      outData_24 <= 0;    
      outData_25 <= 0;    
      outData_26 <= 0;    
      outData_27 <= 0;    
      outData_28 <= 0;    
      outData_29 <= 0;    
      outData_30 <= 0;    
      outData_31 <= 0;    
      outData_32 <= 0;    
      outData_33 <= 0;    
      outData_34 <= 0;    
      outData_35 <= 0;    
      outData_36 <= 0;    
      outData_37 <= 0;    
      outData_38 <= 0;    
      outData_39 <= 0;    
      outData_40 <= 0;    
      outData_41 <= 0;    
      outData_42 <= 0;    
      outData_43 <= 0;    
      outData_44 <= 0;    
      outData_45 <= 0;    
      outData_46 <= 0;    
      outData_47 <= 0;    
      outData_48 <= 0;    
      outData_49 <= 0;    
      outData_50 <= 0;    
      outData_51 <= 0;    
      outData_52 <= 0;    
      outData_53 <= 0;    
      outData_54 <= 0;    
      outData_55 <= 0;    
      outData_56 <= 0;    
      outData_57 <= 0;    
      outData_58 <= 0;    
      outData_59 <= 0;    
      outData_60 <= 0;    
      outData_61 <= 0;    
      outData_62 <= 0;    
      outData_63 <= 0;    
      outData_64 <= 0;    
      outData_65 <= 0;    
      outData_66 <= 0;    
      outData_67 <= 0;    
      outData_68 <= 0;    
      outData_69 <= 0;    
      outData_70 <= 0;    
      outData_71 <= 0;    
      outData_72 <= 0;    
      outData_73 <= 0;    
      outData_74 <= 0;    
      outData_75 <= 0;    
      outData_76 <= 0;    
      outData_77 <= 0;    
      outData_78 <= 0;    
      outData_79 <= 0;    
      outData_80 <= 0;    
      outData_81 <= 0;    
      outData_82 <= 0;    
      outData_83 <= 0;    
      outData_84 <= 0;    
      outData_85 <= 0;    
      outData_86 <= 0;    
      outData_87 <= 0;    
      outData_88 <= 0;    
      outData_89 <= 0;    
      outData_90 <= 0;    
      outData_91 <= 0;    
      outData_92 <= 0;    
      outData_93 <= 0;    
      outData_94 <= 0;    
      outData_95 <= 0;    
      outData_96 <= 0;    
      outData_97 <= 0;    
      outData_98 <= 0;    
      outData_99 <= 0;    
      outData_100 <= 0;    
      outData_101 <= 0;    
      outData_102 <= 0;    
      outData_103 <= 0;    
      outData_104 <= 0;    
      outData_105 <= 0;    
      outData_106 <= 0;    
      outData_107 <= 0;    
      outData_108 <= 0;    
      outData_109 <= 0;    
      outData_110 <= 0;    
      outData_111 <= 0;    
      outData_112 <= 0;    
      outData_113 <= 0;    
      outData_114 <= 0;    
      outData_115 <= 0;    
      outData_116 <= 0;    
      outData_117 <= 0;    
      outData_118 <= 0;    
      outData_119 <= 0;    
      outData_120 <= 0;    
      outData_121 <= 0;    
      outData_122 <= 0;    
      outData_123 <= 0;    
      outData_124 <= 0;    
      outData_125 <= 0;    
      outData_126 <= 0;    
      outData_127 <= 0;    
      outData_128 <= 0;    
      outData_129 <= 0;    
      outData_130 <= 0;    
      outData_131 <= 0;    
      outData_132 <= 0;    
      outData_133 <= 0;    
      outData_134 <= 0;    
      outData_135 <= 0;    
      outData_136 <= 0;    
      outData_137 <= 0;    
      outData_138 <= 0;    
      outData_139 <= 0;    
      outData_140 <= 0;    
      outData_141 <= 0;    
      outData_142 <= 0;    
      outData_143 <= 0;    
      outData_144 <= 0;    
      outData_145 <= 0;    
      outData_146 <= 0;    
      outData_147 <= 0;    
      outData_148 <= 0;    
      outData_149 <= 0;    
      outData_150 <= 0;    
      outData_151 <= 0;    
      outData_152 <= 0;    
      outData_153 <= 0;    
      outData_154 <= 0;    
      outData_155 <= 0;    
      outData_156 <= 0;    
      outData_157 <= 0;    
      outData_158 <= 0;    
      outData_159 <= 0;    
      outData_160 <= 0;    
      outData_161 <= 0;    
      outData_162 <= 0;    
      outData_163 <= 0;    
      outData_164 <= 0;    
      outData_165 <= 0;    
      outData_166 <= 0;    
      outData_167 <= 0;    
      outData_168 <= 0;    
      outData_169 <= 0;    
      outData_170 <= 0;    
      outData_171 <= 0;    
      outData_172 <= 0;    
      outData_173 <= 0;    
      outData_174 <= 0;    
      outData_175 <= 0;    
      outData_176 <= 0;    
      outData_177 <= 0;    
      outData_178 <= 0;    
      outData_179 <= 0;    
      outData_180 <= 0;    
      outData_181 <= 0;    
      outData_182 <= 0;    
      outData_183 <= 0;    
      outData_184 <= 0;    
      outData_185 <= 0;    
      outData_186 <= 0;    
      outData_187 <= 0;    
      outData_188 <= 0;    
      outData_189 <= 0;    
      outData_190 <= 0;    
      outData_191 <= 0;    
      outData_192 <= 0;    
      outData_193 <= 0;    
      outData_194 <= 0;    
      outData_195 <= 0;    
      outData_196 <= 0;    
      outData_197 <= 0;    
      outData_198 <= 0;    
      outData_199 <= 0;    
      outData_200 <= 0;    
      outData_201 <= 0;    
      outData_202 <= 0;    
      outData_203 <= 0;    
      outData_204 <= 0;    
      outData_205 <= 0;    
      outData_206 <= 0;    
      outData_207 <= 0;    
      outData_208 <= 0;    
      outData_209 <= 0;    
      outData_210 <= 0;    
      outData_211 <= 0;    
      outData_212 <= 0;    
      outData_213 <= 0;    
      outData_214 <= 0;    
      outData_215 <= 0;    
      outData_216 <= 0;    
      outData_217 <= 0;    
      outData_218 <= 0;    
      outData_219 <= 0;    
      outData_220 <= 0;    
      outData_221 <= 0;    
      outData_222 <= 0;    
      outData_223 <= 0;    
      outData_224 <= 0;    
      outData_225 <= 0;    
      outData_226 <= 0;    
      outData_227 <= 0;    
      outData_228 <= 0;    
      outData_229 <= 0;    
      outData_230 <= 0;    
      outData_231 <= 0;    
      outData_232 <= 0;    
      outData_233 <= 0;    
      outData_234 <= 0;    
      outData_235 <= 0;    
      outData_236 <= 0;    
      outData_237 <= 0;    
      outData_238 <= 0;    
      outData_239 <= 0;    
      outData_240 <= 0;    
      outData_241 <= 0;    
      outData_242 <= 0;    
      outData_243 <= 0;    
      outData_244 <= 0;    
      outData_245 <= 0;    
      outData_246 <= 0;    
      outData_247 <= 0;    
      outData_248 <= 0;    
      outData_249 <= 0;    
      outData_250 <= 0;    
      outData_251 <= 0;    
      outData_252 <= 0;    
      outData_253 <= 0;    
      outData_254 <= 0;    
      outData_255 <= 0;    
      out_start <= 1'b0;    
      end
    else begin                        
      outData_0 <= wireOut[0];    
      outData_1 <= wireOut[1];    
      outData_2 <= wireOut[2];    
      outData_3 <= wireOut[3];    
      outData_4 <= wireOut[4];    
      outData_5 <= wireOut[5];    
      outData_6 <= wireOut[6];    
      outData_7 <= wireOut[7];    
      outData_8 <= wireOut[8];    
      outData_9 <= wireOut[9];    
      outData_10 <= wireOut[10];    
      outData_11 <= wireOut[11];    
      outData_12 <= wireOut[12];    
      outData_13 <= wireOut[13];    
      outData_14 <= wireOut[14];    
      outData_15 <= wireOut[15];    
      outData_16 <= wireOut[16];    
      outData_17 <= wireOut[17];    
      outData_18 <= wireOut[18];    
      outData_19 <= wireOut[19];    
      outData_20 <= wireOut[20];    
      outData_21 <= wireOut[21];    
      outData_22 <= wireOut[22];    
      outData_23 <= wireOut[23];    
      outData_24 <= wireOut[24];    
      outData_25 <= wireOut[25];    
      outData_26 <= wireOut[26];    
      outData_27 <= wireOut[27];    
      outData_28 <= wireOut[28];    
      outData_29 <= wireOut[29];    
      outData_30 <= wireOut[30];    
      outData_31 <= wireOut[31];    
      outData_32 <= wireOut[32];    
      outData_33 <= wireOut[33];    
      outData_34 <= wireOut[34];    
      outData_35 <= wireOut[35];    
      outData_36 <= wireOut[36];    
      outData_37 <= wireOut[37];    
      outData_38 <= wireOut[38];    
      outData_39 <= wireOut[39];    
      outData_40 <= wireOut[40];    
      outData_41 <= wireOut[41];    
      outData_42 <= wireOut[42];    
      outData_43 <= wireOut[43];    
      outData_44 <= wireOut[44];    
      outData_45 <= wireOut[45];    
      outData_46 <= wireOut[46];    
      outData_47 <= wireOut[47];    
      outData_48 <= wireOut[48];    
      outData_49 <= wireOut[49];    
      outData_50 <= wireOut[50];    
      outData_51 <= wireOut[51];    
      outData_52 <= wireOut[52];    
      outData_53 <= wireOut[53];    
      outData_54 <= wireOut[54];    
      outData_55 <= wireOut[55];    
      outData_56 <= wireOut[56];    
      outData_57 <= wireOut[57];    
      outData_58 <= wireOut[58];    
      outData_59 <= wireOut[59];    
      outData_60 <= wireOut[60];    
      outData_61 <= wireOut[61];    
      outData_62 <= wireOut[62];    
      outData_63 <= wireOut[63];    
      outData_64 <= wireOut[64];    
      outData_65 <= wireOut[65];    
      outData_66 <= wireOut[66];    
      outData_67 <= wireOut[67];    
      outData_68 <= wireOut[68];    
      outData_69 <= wireOut[69];    
      outData_70 <= wireOut[70];    
      outData_71 <= wireOut[71];    
      outData_72 <= wireOut[72];    
      outData_73 <= wireOut[73];    
      outData_74 <= wireOut[74];    
      outData_75 <= wireOut[75];    
      outData_76 <= wireOut[76];    
      outData_77 <= wireOut[77];    
      outData_78 <= wireOut[78];    
      outData_79 <= wireOut[79];    
      outData_80 <= wireOut[80];    
      outData_81 <= wireOut[81];    
      outData_82 <= wireOut[82];    
      outData_83 <= wireOut[83];    
      outData_84 <= wireOut[84];    
      outData_85 <= wireOut[85];    
      outData_86 <= wireOut[86];    
      outData_87 <= wireOut[87];    
      outData_88 <= wireOut[88];    
      outData_89 <= wireOut[89];    
      outData_90 <= wireOut[90];    
      outData_91 <= wireOut[91];    
      outData_92 <= wireOut[92];    
      outData_93 <= wireOut[93];    
      outData_94 <= wireOut[94];    
      outData_95 <= wireOut[95];    
      outData_96 <= wireOut[96];    
      outData_97 <= wireOut[97];    
      outData_98 <= wireOut[98];    
      outData_99 <= wireOut[99];    
      outData_100 <= wireOut[100];    
      outData_101 <= wireOut[101];    
      outData_102 <= wireOut[102];    
      outData_103 <= wireOut[103];    
      outData_104 <= wireOut[104];    
      outData_105 <= wireOut[105];    
      outData_106 <= wireOut[106];    
      outData_107 <= wireOut[107];    
      outData_108 <= wireOut[108];    
      outData_109 <= wireOut[109];    
      outData_110 <= wireOut[110];    
      outData_111 <= wireOut[111];    
      outData_112 <= wireOut[112];    
      outData_113 <= wireOut[113];    
      outData_114 <= wireOut[114];    
      outData_115 <= wireOut[115];    
      outData_116 <= wireOut[116];    
      outData_117 <= wireOut[117];    
      outData_118 <= wireOut[118];    
      outData_119 <= wireOut[119];    
      outData_120 <= wireOut[120];    
      outData_121 <= wireOut[121];    
      outData_122 <= wireOut[122];    
      outData_123 <= wireOut[123];    
      outData_124 <= wireOut[124];    
      outData_125 <= wireOut[125];    
      outData_126 <= wireOut[126];    
      outData_127 <= wireOut[127];    
      outData_128 <= wireOut[128];    
      outData_129 <= wireOut[129];    
      outData_130 <= wireOut[130];    
      outData_131 <= wireOut[131];    
      outData_132 <= wireOut[132];    
      outData_133 <= wireOut[133];    
      outData_134 <= wireOut[134];    
      outData_135 <= wireOut[135];    
      outData_136 <= wireOut[136];    
      outData_137 <= wireOut[137];    
      outData_138 <= wireOut[138];    
      outData_139 <= wireOut[139];    
      outData_140 <= wireOut[140];    
      outData_141 <= wireOut[141];    
      outData_142 <= wireOut[142];    
      outData_143 <= wireOut[143];    
      outData_144 <= wireOut[144];    
      outData_145 <= wireOut[145];    
      outData_146 <= wireOut[146];    
      outData_147 <= wireOut[147];    
      outData_148 <= wireOut[148];    
      outData_149 <= wireOut[149];    
      outData_150 <= wireOut[150];    
      outData_151 <= wireOut[151];    
      outData_152 <= wireOut[152];    
      outData_153 <= wireOut[153];    
      outData_154 <= wireOut[154];    
      outData_155 <= wireOut[155];    
      outData_156 <= wireOut[156];    
      outData_157 <= wireOut[157];    
      outData_158 <= wireOut[158];    
      outData_159 <= wireOut[159];    
      outData_160 <= wireOut[160];    
      outData_161 <= wireOut[161];    
      outData_162 <= wireOut[162];    
      outData_163 <= wireOut[163];    
      outData_164 <= wireOut[164];    
      outData_165 <= wireOut[165];    
      outData_166 <= wireOut[166];    
      outData_167 <= wireOut[167];    
      outData_168 <= wireOut[168];    
      outData_169 <= wireOut[169];    
      outData_170 <= wireOut[170];    
      outData_171 <= wireOut[171];    
      outData_172 <= wireOut[172];    
      outData_173 <= wireOut[173];    
      outData_174 <= wireOut[174];    
      outData_175 <= wireOut[175];    
      outData_176 <= wireOut[176];    
      outData_177 <= wireOut[177];    
      outData_178 <= wireOut[178];    
      outData_179 <= wireOut[179];    
      outData_180 <= wireOut[180];    
      outData_181 <= wireOut[181];    
      outData_182 <= wireOut[182];    
      outData_183 <= wireOut[183];    
      outData_184 <= wireOut[184];    
      outData_185 <= wireOut[185];    
      outData_186 <= wireOut[186];    
      outData_187 <= wireOut[187];    
      outData_188 <= wireOut[188];    
      outData_189 <= wireOut[189];    
      outData_190 <= wireOut[190];    
      outData_191 <= wireOut[191];    
      outData_192 <= wireOut[192];    
      outData_193 <= wireOut[193];    
      outData_194 <= wireOut[194];    
      outData_195 <= wireOut[195];    
      outData_196 <= wireOut[196];    
      outData_197 <= wireOut[197];    
      outData_198 <= wireOut[198];    
      outData_199 <= wireOut[199];    
      outData_200 <= wireOut[200];    
      outData_201 <= wireOut[201];    
      outData_202 <= wireOut[202];    
      outData_203 <= wireOut[203];    
      outData_204 <= wireOut[204];    
      outData_205 <= wireOut[205];    
      outData_206 <= wireOut[206];    
      outData_207 <= wireOut[207];    
      outData_208 <= wireOut[208];    
      outData_209 <= wireOut[209];    
      outData_210 <= wireOut[210];    
      outData_211 <= wireOut[211];    
      outData_212 <= wireOut[212];    
      outData_213 <= wireOut[213];    
      outData_214 <= wireOut[214];    
      outData_215 <= wireOut[215];    
      outData_216 <= wireOut[216];    
      outData_217 <= wireOut[217];    
      outData_218 <= wireOut[218];    
      outData_219 <= wireOut[219];    
      outData_220 <= wireOut[220];    
      outData_221 <= wireOut[221];    
      outData_222 <= wireOut[222];    
      outData_223 <= wireOut[223];    
      outData_224 <= wireOut[224];    
      outData_225 <= wireOut[225];    
      outData_226 <= wireOut[226];    
      outData_227 <= wireOut[227];    
      outData_228 <= wireOut[228];    
      outData_229 <= wireOut[229];    
      outData_230 <= wireOut[230];    
      outData_231 <= wireOut[231];    
      outData_232 <= wireOut[232];    
      outData_233 <= wireOut[233];    
      outData_234 <= wireOut[234];    
      outData_235 <= wireOut[235];    
      outData_236 <= wireOut[236];    
      outData_237 <= wireOut[237];    
      outData_238 <= wireOut[238];    
      outData_239 <= wireOut[239];    
      outData_240 <= wireOut[240];    
      outData_241 <= wireOut[241];    
      outData_242 <= wireOut[242];    
      outData_243 <= wireOut[243];    
      outData_244 <= wireOut[244];    
      outData_245 <= wireOut[245];    
      outData_246 <= wireOut[246];    
      outData_247 <= wireOut[247];    
      outData_248 <= wireOut[248];    
      outData_249 <= wireOut[249];    
      outData_250 <= wireOut[250];    
      outData_251 <= wireOut[251];    
      outData_252 <= wireOut[252];    
      outData_253 <= wireOut[253];    
      outData_254 <= wireOut[254];    
      outData_255 <= wireOut[255];    
      out_start <= out_start_RB;    
      end
  end                              

endmodule                        

